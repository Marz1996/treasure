
module mR4000 ( Clk, Reset, MemData, ReadAdd, WriteAdd, WriteData, MemWrite, 
        MemRead );
  input [31:0] MemData;
  output [31:0] ReadAdd;
  output [31:0] WriteAdd;
  output [31:0] WriteData;
  input Clk, Reset;
  output MemWrite, MemRead;
  wire   Instruction_31, Instruction_30, Instruction_29, Instruction_28,
         Instruction_27, Instruction_26, Instruction_25, Instruction_24,
         Instruction_23, Instruction_20, Instruction_19, Instruction_18,
         RegDst, MemToReg, IRWrite, PCWriteCond, PCWrite, TargetWrite, IorD,
         RegWrite, cntrl_N116, cntrl_N114, cntrl_N113, cntrl_N111, cntrl_N109,
         cntrl_N106, cntrl_N104, cntrl_N103, cntrl_state_0_, cntrl_state_1_,
         cntrl_state_2_, cntrl_state_3_, cntrl_state_4_, cntrl_state_5_,
         cntrl_state_6_, cntrl_state_7_, cntrl_state_8_, cntrl_state_9_,
         cntrl_state_10_, alu_MuxB_1_, alu_MuxB_2_, alu_MuxB_3_, alu_MuxB_4_,
         alu_MuxB_5_, alu_MuxB_6_, alu_MuxB_7_, alu_MuxB_8_, alu_MuxB_9_,
         alu_MuxB_10_, alu_MuxB_11_, alu_MuxB_12_, alu_MuxB_13_, alu_MuxB_14_,
         alu_MuxB_15_, alu_MuxB_16_, alu_MuxB_17_, alu_MuxB_18_, alu_MuxB_19_,
         alu_MuxB_20_, alu_MuxB_21_, alu_MuxB_22_, alu_MuxB_23_, alu_MuxB_24_,
         alu_MuxB_25_, alu_MuxB_26_, alu_MuxB_27_, alu_MuxB_28_, alu_MuxB_29_,
         alu_MuxB_30_, alu_MuxB_31_, alu_MuxA_0_, alu_MuxA_1_, alu_MuxA_2_,
         alu_MuxA_3_, alu_MuxA_4_, alu_MuxA_5_, alu_MuxA_6_, alu_MuxA_7_,
         alu_MuxA_8_, alu_MuxA_9_, alu_MuxA_10_, alu_MuxA_11_, alu_MuxA_12_,
         alu_MuxA_13_, alu_MuxA_14_, alu_MuxA_15_, alu_MuxA_16_, alu_MuxA_17_,
         alu_MuxA_18_, alu_MuxA_19_, alu_MuxA_20_, alu_MuxA_21_, alu_MuxA_22_,
         alu_MuxA_23_, alu_MuxA_24_, alu_MuxA_25_, alu_MuxA_26_, alu_MuxA_27_,
         alu_MuxA_28_, alu_MuxA_29_, alu_MuxA_30_, alu_MuxA_31_, C55_DATA6_0,
         C55_DATA6_1, C55_DATA6_2, C55_DATA6_3, C55_DATA6_4, C55_DATA6_5,
         C55_DATA6_6, C55_DATA6_7, C55_DATA6_8, C55_DATA6_9, C55_DATA6_10,
         C55_DATA6_11, C55_DATA6_12, C55_DATA6_13, C55_DATA6_14, C55_DATA6_15,
         C55_DATA6_16, C55_DATA6_17, C55_DATA6_18, C55_DATA6_19, C55_DATA6_20,
         C55_DATA6_21, C55_DATA6_22, C55_DATA6_23, C55_DATA6_24, C55_DATA6_25,
         C55_DATA6_26, C55_DATA6_27, C55_DATA6_28, C55_DATA6_29, C55_DATA6_30,
         C55_DATA6_31, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n139, n140, n142,
         n144, n145, n155, n156, n157, n419, n426, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, DP_OP_100J1_124_3689_n100,
         DP_OP_100J1_124_3689_n66, DP_OP_100J1_124_3689_n65,
         DP_OP_100J1_124_3689_n64, DP_OP_100J1_124_3689_n63,
         DP_OP_100J1_124_3689_n62, DP_OP_100J1_124_3689_n61,
         DP_OP_100J1_124_3689_n60, DP_OP_100J1_124_3689_n59,
         DP_OP_100J1_124_3689_n58, DP_OP_100J1_124_3689_n57,
         DP_OP_100J1_124_3689_n56, DP_OP_100J1_124_3689_n55,
         DP_OP_100J1_124_3689_n54, DP_OP_100J1_124_3689_n53,
         DP_OP_100J1_124_3689_n52, DP_OP_100J1_124_3689_n51,
         DP_OP_100J1_124_3689_n50, DP_OP_100J1_124_3689_n49,
         DP_OP_100J1_124_3689_n48, DP_OP_100J1_124_3689_n47,
         DP_OP_100J1_124_3689_n46, DP_OP_100J1_124_3689_n45,
         DP_OP_100J1_124_3689_n44, DP_OP_100J1_124_3689_n43,
         DP_OP_100J1_124_3689_n42, DP_OP_100J1_124_3689_n41,
         DP_OP_100J1_124_3689_n40, DP_OP_100J1_124_3689_n39,
         DP_OP_100J1_124_3689_n38, DP_OP_100J1_124_3689_n37,
         DP_OP_100J1_124_3689_n36, DP_OP_100J1_124_3689_n31,
         DP_OP_100J1_124_3689_n30, DP_OP_100J1_124_3689_n29,
         DP_OP_100J1_124_3689_n28, DP_OP_100J1_124_3689_n27,
         DP_OP_100J1_124_3689_n26, DP_OP_100J1_124_3689_n25,
         DP_OP_100J1_124_3689_n24, DP_OP_100J1_124_3689_n23,
         DP_OP_100J1_124_3689_n22, DP_OP_100J1_124_3689_n21,
         DP_OP_100J1_124_3689_n20, DP_OP_100J1_124_3689_n19,
         DP_OP_100J1_124_3689_n18, DP_OP_100J1_124_3689_n17,
         DP_OP_100J1_124_3689_n16, DP_OP_100J1_124_3689_n15,
         DP_OP_100J1_124_3689_n14, DP_OP_100J1_124_3689_n13,
         DP_OP_100J1_124_3689_n12, DP_OP_100J1_124_3689_n11,
         DP_OP_100J1_124_3689_n10, DP_OP_100J1_124_3689_n9,
         DP_OP_100J1_124_3689_n8, DP_OP_100J1_124_3689_n7,
         DP_OP_100J1_124_3689_n6, DP_OP_100J1_124_3689_n5,
         DP_OP_100J1_124_3689_n4, DP_OP_100J1_124_3689_n3,
         DP_OP_100J1_124_3689_n2, DP_OP_100J1_124_3689_n1, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481;
  wire   [1:0] Read1RegSel;
  wire   [15:0] Instruction;
  wire   [1:0] Read2RegSel;
  wire   [1:0] PCSource;
  wire   [31:0] PC;
  wire   [31:0] TargetReg;
  wire   [1:0] ALUOp;
  wire   [1:0] ALUSelB;

  fa1b0 DP_OP_100J1_124_3689_U31 ( .CI(DP_OP_100J1_124_3689_n31), .B(
        alu_MuxA_1_), .A(DP_OP_100J1_124_3689_n66), .S(C55_DATA6_1), .CO(
        DP_OP_100J1_124_3689_n30) );
  fa2a0 DP_OP_100J1_124_3689_U30 ( .A(DP_OP_100J1_124_3689_n65), .B(
        alu_MuxA_2_), .CI(DP_OP_100J1_124_3689_n30), .CO(
        DP_OP_100J1_124_3689_n29), .S(C55_DATA6_2) );
  fa1b0 DP_OP_100J1_124_3689_U29 ( .CI(DP_OP_100J1_124_3689_n29), .B(
        alu_MuxA_3_), .A(DP_OP_100J1_124_3689_n64), .S(C55_DATA6_3), .CO(
        DP_OP_100J1_124_3689_n28) );
  fa2a0 DP_OP_100J1_124_3689_U28 ( .A(DP_OP_100J1_124_3689_n63), .B(
        alu_MuxA_4_), .CI(DP_OP_100J1_124_3689_n28), .CO(
        DP_OP_100J1_124_3689_n27), .S(C55_DATA6_4) );
  fa1b0 DP_OP_100J1_124_3689_U27 ( .CI(DP_OP_100J1_124_3689_n27), .B(
        alu_MuxA_5_), .A(DP_OP_100J1_124_3689_n62), .S(C55_DATA6_5), .CO(
        DP_OP_100J1_124_3689_n26) );
  fa2a0 DP_OP_100J1_124_3689_U26 ( .A(DP_OP_100J1_124_3689_n61), .B(
        alu_MuxA_6_), .CI(DP_OP_100J1_124_3689_n26), .CO(
        DP_OP_100J1_124_3689_n25), .S(C55_DATA6_6) );
  fa1b0 DP_OP_100J1_124_3689_U25 ( .CI(DP_OP_100J1_124_3689_n25), .B(
        alu_MuxA_7_), .A(DP_OP_100J1_124_3689_n60), .S(C55_DATA6_7), .CO(
        DP_OP_100J1_124_3689_n24) );
  fa2a0 DP_OP_100J1_124_3689_U24 ( .A(DP_OP_100J1_124_3689_n59), .B(
        alu_MuxA_8_), .CI(DP_OP_100J1_124_3689_n24), .CO(
        DP_OP_100J1_124_3689_n23), .S(C55_DATA6_8) );
  fa1b0 DP_OP_100J1_124_3689_U23 ( .CI(DP_OP_100J1_124_3689_n23), .B(
        alu_MuxA_9_), .A(DP_OP_100J1_124_3689_n58), .S(C55_DATA6_9), .CO(
        DP_OP_100J1_124_3689_n22) );
  fa2a0 DP_OP_100J1_124_3689_U22 ( .A(DP_OP_100J1_124_3689_n57), .B(
        alu_MuxA_10_), .CI(DP_OP_100J1_124_3689_n22), .CO(
        DP_OP_100J1_124_3689_n21), .S(C55_DATA6_10) );
  fa1b0 DP_OP_100J1_124_3689_U21 ( .CI(DP_OP_100J1_124_3689_n21), .B(
        alu_MuxA_11_), .A(DP_OP_100J1_124_3689_n56), .S(C55_DATA6_11), .CO(
        DP_OP_100J1_124_3689_n20) );
  fa2a0 DP_OP_100J1_124_3689_U20 ( .A(DP_OP_100J1_124_3689_n55), .B(
        alu_MuxA_12_), .CI(DP_OP_100J1_124_3689_n20), .CO(
        DP_OP_100J1_124_3689_n19), .S(C55_DATA6_12) );
  fa1b0 DP_OP_100J1_124_3689_U19 ( .CI(DP_OP_100J1_124_3689_n19), .B(
        alu_MuxA_13_), .A(DP_OP_100J1_124_3689_n54), .S(C55_DATA6_13), .CO(
        DP_OP_100J1_124_3689_n18) );
  fa2a0 DP_OP_100J1_124_3689_U18 ( .A(DP_OP_100J1_124_3689_n53), .B(
        alu_MuxA_14_), .CI(DP_OP_100J1_124_3689_n18), .CO(
        DP_OP_100J1_124_3689_n17), .S(C55_DATA6_14) );
  fa1b0 DP_OP_100J1_124_3689_U17 ( .CI(DP_OP_100J1_124_3689_n17), .B(
        alu_MuxA_15_), .A(DP_OP_100J1_124_3689_n52), .S(C55_DATA6_15), .CO(
        DP_OP_100J1_124_3689_n16) );
  fa2a0 DP_OP_100J1_124_3689_U16 ( .A(DP_OP_100J1_124_3689_n51), .B(
        alu_MuxA_16_), .CI(DP_OP_100J1_124_3689_n16), .CO(
        DP_OP_100J1_124_3689_n15), .S(C55_DATA6_16) );
  fa1b0 DP_OP_100J1_124_3689_U15 ( .CI(DP_OP_100J1_124_3689_n15), .B(
        alu_MuxA_17_), .A(DP_OP_100J1_124_3689_n50), .S(C55_DATA6_17), .CO(
        DP_OP_100J1_124_3689_n14) );
  fa2a0 DP_OP_100J1_124_3689_U14 ( .A(DP_OP_100J1_124_3689_n49), .B(
        alu_MuxA_18_), .CI(DP_OP_100J1_124_3689_n14), .CO(
        DP_OP_100J1_124_3689_n13), .S(C55_DATA6_18) );
  fa1b0 DP_OP_100J1_124_3689_U13 ( .CI(DP_OP_100J1_124_3689_n13), .B(
        alu_MuxA_19_), .A(DP_OP_100J1_124_3689_n48), .S(C55_DATA6_19), .CO(
        DP_OP_100J1_124_3689_n12) );
  fa2a0 DP_OP_100J1_124_3689_U12 ( .A(DP_OP_100J1_124_3689_n47), .B(
        alu_MuxA_20_), .CI(DP_OP_100J1_124_3689_n12), .CO(
        DP_OP_100J1_124_3689_n11), .S(C55_DATA6_20) );
  fa1b0 DP_OP_100J1_124_3689_U11 ( .CI(DP_OP_100J1_124_3689_n11), .B(
        alu_MuxA_21_), .A(DP_OP_100J1_124_3689_n46), .S(C55_DATA6_21), .CO(
        DP_OP_100J1_124_3689_n10) );
  fa2a0 DP_OP_100J1_124_3689_U10 ( .A(DP_OP_100J1_124_3689_n45), .B(
        alu_MuxA_22_), .CI(DP_OP_100J1_124_3689_n10), .CO(
        DP_OP_100J1_124_3689_n9), .S(C55_DATA6_22) );
  fa1b0 DP_OP_100J1_124_3689_U9 ( .CI(DP_OP_100J1_124_3689_n9), .B(
        alu_MuxA_23_), .A(DP_OP_100J1_124_3689_n44), .S(C55_DATA6_23), .CO(
        DP_OP_100J1_124_3689_n8) );
  fa2a0 DP_OP_100J1_124_3689_U8 ( .A(DP_OP_100J1_124_3689_n43), .B(
        alu_MuxA_24_), .CI(DP_OP_100J1_124_3689_n8), .CO(
        DP_OP_100J1_124_3689_n7), .S(C55_DATA6_24) );
  fa1b0 DP_OP_100J1_124_3689_U7 ( .CI(DP_OP_100J1_124_3689_n7), .B(
        alu_MuxA_25_), .A(DP_OP_100J1_124_3689_n42), .S(C55_DATA6_25), .CO(
        DP_OP_100J1_124_3689_n6) );
  fa2a0 DP_OP_100J1_124_3689_U6 ( .A(DP_OP_100J1_124_3689_n41), .B(
        alu_MuxA_26_), .CI(DP_OP_100J1_124_3689_n6), .CO(
        DP_OP_100J1_124_3689_n5), .S(C55_DATA6_26) );
  fa1b0 DP_OP_100J1_124_3689_U5 ( .CI(DP_OP_100J1_124_3689_n5), .B(
        alu_MuxA_27_), .A(DP_OP_100J1_124_3689_n40), .S(C55_DATA6_27), .CO(
        DP_OP_100J1_124_3689_n4) );
  fa2a0 DP_OP_100J1_124_3689_U4 ( .A(DP_OP_100J1_124_3689_n39), .B(
        alu_MuxA_28_), .CI(DP_OP_100J1_124_3689_n4), .CO(
        DP_OP_100J1_124_3689_n3), .S(C55_DATA6_28) );
  fa1b0 DP_OP_100J1_124_3689_U3 ( .CI(DP_OP_100J1_124_3689_n3), .B(
        alu_MuxA_29_), .A(DP_OP_100J1_124_3689_n38), .S(C55_DATA6_29), .CO(
        DP_OP_100J1_124_3689_n2) );
  fa2a0 DP_OP_100J1_124_3689_U2 ( .A(DP_OP_100J1_124_3689_n37), .B(
        alu_MuxA_30_), .CI(DP_OP_100J1_124_3689_n2), .CO(
        DP_OP_100J1_124_3689_n1), .S(C55_DATA6_30) );
  fa1b0 DP_OP_100J1_124_3689_U1 ( .CI(DP_OP_100J1_124_3689_n1), .B(
        alu_MuxA_31_), .A(DP_OP_100J1_124_3689_n36), .S(C55_DATA6_31) );
  fdm5a2 cntrl_IorD_reg ( .D0(cntrl_state_2_), .D1(n144), .D2(n142), .S0(
        cntrl_state_1_), .S1(Reset), .CLK(Clk), .Q(IorD) );
  fd1c2 cntrl_ALUSelA_reg ( .D(cntrl_N113), .CLK(Clk), .QN(n139) );
  fd1a2 cntrl_TargetWrite_reg ( .D(cntrl_N116), .CLK(Clk), .Q(TargetWrite) );
  fdm5a2 cntrl_IRWrite_reg ( .D0(cntrl_state_7_), .D1(n144), .D2(n144), .S0(
        n426), .S1(Reset), .CLK(Clk), .Q(IRWrite) );
  fd1a2 cntrl_MemWrite_reg ( .D(cntrl_N103), .CLK(Clk), .Q(MemWrite) );
  fd1a2 cntrl_MemRead_reg ( .D(cntrl_N104), .CLK(Clk), .Q(MemRead) );
  fd1a2 cntrl_state_reg_4_ ( .D(n897), .CLK(Clk), .Q(cntrl_state_4_) );
  fd1a2 cntrl_state_reg_5_ ( .D(cntrl_N103), .CLK(Clk), .Q(cntrl_state_5_) );
  fd1a2 cntrl_PCWriteCond_reg ( .D(cntrl_N106), .CLK(Clk), .Q(PCWriteCond) );
  fdm5a2 cntrl_PCWrite_reg ( .D0(n142), .D1(n971), .D2(n144), .S0(
        cntrl_state_0_), .S1(n900), .CLK(Clk), .Q(PCWrite) );
  fde1a2 Instruction_reg_18_ ( .D(MemData[18]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction_18) );
  fde1a2 Instruction_reg_19_ ( .D(MemData[19]), .E(n978), .CLK(Clk), .Q(
        Instruction_19) );
  fde1a2 Instruction_reg_20_ ( .D(MemData[20]), .E(n977), .CLK(Clk), .Q(
        Instruction_20) );
  fde1a2 Instruction_reg_23_ ( .D(MemData[23]), .E(n978), .CLK(Clk), .Q(
        Instruction_23) );
  fde1a2 Instruction_reg_24_ ( .D(MemData[24]), .E(n977), .CLK(Clk), .Q(
        Instruction_24) );
  fde1a2 Instruction_reg_25_ ( .D(MemData[25]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction_25) );
  fde1a2 TargetReg_reg_2_ ( .D(WriteAdd[2]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[2]) );
  fde1a2 TargetReg_reg_1_ ( .D(WriteAdd[1]), .E(n976), .CLK(Clk), .Q(
        TargetReg[1]) );
  fde1a2 TargetReg_reg_0_ ( .D(WriteAdd[0]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[0]) );
  fde1a2 TargetReg_reg_31_ ( .D(WriteAdd[31]), .E(n976), .CLK(Clk), .Q(
        TargetReg[31]) );
  fde1a2 TargetReg_reg_30_ ( .D(WriteAdd[30]), .E(n975), .CLK(Clk), .Q(
        TargetReg[30]) );
  fde1a2 TargetReg_reg_27_ ( .D(WriteAdd[27]), .E(n976), .CLK(Clk), .Q(
        TargetReg[27]) );
  fde1a2 TargetReg_reg_28_ ( .D(WriteAdd[28]), .E(n976), .CLK(Clk), .Q(
        TargetReg[28]) );
  fde1a2 TargetReg_reg_29_ ( .D(WriteAdd[29]), .E(n976), .CLK(Clk), .Q(
        TargetReg[29]) );
  fde1a2 TargetReg_reg_26_ ( .D(WriteAdd[26]), .E(n975), .CLK(Clk), .Q(
        TargetReg[26]) );
  fde1a2 TargetReg_reg_25_ ( .D(WriteAdd[25]), .E(n975), .CLK(Clk), .Q(
        TargetReg[25]) );
  fde1a2 TargetReg_reg_24_ ( .D(WriteAdd[24]), .E(n975), .CLK(Clk), .Q(
        TargetReg[24]) );
  fde1a2 TargetReg_reg_23_ ( .D(WriteAdd[23]), .E(n975), .CLK(Clk), .Q(
        TargetReg[23]) );
  fde1a2 TargetReg_reg_22_ ( .D(WriteAdd[22]), .E(n975), .CLK(Clk), .Q(
        TargetReg[22]) );
  fde1a2 TargetReg_reg_21_ ( .D(WriteAdd[21]), .E(n975), .CLK(Clk), .Q(
        TargetReg[21]) );
  fde1a2 TargetReg_reg_20_ ( .D(WriteAdd[20]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[20]) );
  fde1a2 TargetReg_reg_19_ ( .D(WriteAdd[19]), .E(n976), .CLK(Clk), .Q(
        TargetReg[19]) );
  fde1a2 TargetReg_reg_18_ ( .D(WriteAdd[18]), .E(n975), .CLK(Clk), .Q(
        TargetReg[18]) );
  fde1a2 TargetReg_reg_17_ ( .D(WriteAdd[17]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[17]) );
  fde1a2 TargetReg_reg_16_ ( .D(WriteAdd[16]), .E(n976), .CLK(Clk), .Q(
        TargetReg[16]) );
  fde1a2 TargetReg_reg_15_ ( .D(WriteAdd[15]), .E(n975), .CLK(Clk), .Q(
        TargetReg[15]) );
  fde1a2 TargetReg_reg_14_ ( .D(WriteAdd[14]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[14]) );
  fde1a2 TargetReg_reg_13_ ( .D(WriteAdd[13]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[13]) );
  fde1a2 TargetReg_reg_12_ ( .D(WriteAdd[12]), .E(n976), .CLK(Clk), .Q(
        TargetReg[12]) );
  fde1a2 TargetReg_reg_11_ ( .D(WriteAdd[11]), .E(n975), .CLK(Clk), .Q(
        TargetReg[11]) );
  fde1a2 TargetReg_reg_10_ ( .D(WriteAdd[10]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[10]) );
  fde1a2 TargetReg_reg_9_ ( .D(WriteAdd[9]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[9]) );
  fde1a2 TargetReg_reg_8_ ( .D(WriteAdd[8]), .E(n976), .CLK(Clk), .Q(
        TargetReg[8]) );
  fde1a2 TargetReg_reg_7_ ( .D(WriteAdd[7]), .E(n975), .CLK(Clk), .Q(
        TargetReg[7]) );
  fde1a2 TargetReg_reg_6_ ( .D(WriteAdd[6]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[6]) );
  fde1a2 TargetReg_reg_5_ ( .D(WriteAdd[5]), .E(n976), .CLK(Clk), .Q(
        TargetReg[5]) );
  fde1a2 TargetReg_reg_4_ ( .D(WriteAdd[4]), .E(TargetWrite), .CLK(Clk), .Q(
        TargetReg[4]) );
  fde1a2 TargetReg_reg_3_ ( .D(WriteAdd[3]), .E(n976), .CLK(Clk), .Q(
        TargetReg[3]) );
  fd1c2 register_register1_reg_31_ ( .D(n737), .CLK(Clk), .QN(n126) );
  fd1c2 register_register1_reg_27_ ( .D(n753), .CLK(Clk), .QN(n122) );
  fd1c2 register_register1_reg_28_ ( .D(n749), .CLK(Clk), .QN(n118) );
  fd1c2 register_register1_reg_29_ ( .D(n745), .CLK(Clk), .QN(n114) );
  fd1c2 register_register1_reg_26_ ( .D(n757), .CLK(Clk), .QN(n110) );
  fd1c2 register_register1_reg_25_ ( .D(n761), .CLK(Clk), .QN(n106) );
  fd1c2 register_register1_reg_24_ ( .D(n765), .CLK(Clk), .QN(n102) );
  fd1c2 register_register1_reg_23_ ( .D(n769), .CLK(Clk), .QN(n98) );
  fd1c2 register_register1_reg_22_ ( .D(n773), .CLK(Clk), .QN(n94) );
  fd1c2 register_register1_reg_21_ ( .D(n777), .CLK(Clk), .QN(n90) );
  fd1c2 register_register1_reg_20_ ( .D(n781), .CLK(Clk), .QN(n86) );
  fd1c2 register_register1_reg_19_ ( .D(n785), .CLK(Clk), .QN(n82) );
  fd1c2 register_register1_reg_18_ ( .D(n789), .CLK(Clk), .QN(n78) );
  fd1c2 register_register1_reg_17_ ( .D(n793), .CLK(Clk), .QN(n74) );
  fd1c2 register_register1_reg_16_ ( .D(n797), .CLK(Clk), .QN(n70) );
  fd1c2 register_register1_reg_15_ ( .D(n801), .CLK(Clk), .QN(n66) );
  fd1c2 register_register1_reg_14_ ( .D(n805), .CLK(Clk), .QN(n62) );
  fd1c2 register_register1_reg_13_ ( .D(n809), .CLK(Clk), .QN(n58) );
  fd1c2 register_register1_reg_12_ ( .D(n813), .CLK(Clk), .QN(n54) );
  fd1c2 register_register1_reg_11_ ( .D(n817), .CLK(Clk), .QN(n50) );
  fd1c2 register_register1_reg_10_ ( .D(n821), .CLK(Clk), .QN(n46) );
  fd1c2 register_register1_reg_9_ ( .D(n825), .CLK(Clk), .QN(n42) );
  fd1c2 register_register1_reg_8_ ( .D(n829), .CLK(Clk), .QN(n38) );
  fd1c2 register_register1_reg_7_ ( .D(n833), .CLK(Clk), .QN(n34) );
  fd1c2 register_register1_reg_6_ ( .D(n837), .CLK(Clk), .QN(n30) );
  fd1c2 register_register1_reg_5_ ( .D(n841), .CLK(Clk), .QN(n26) );
  fd1c2 register_register1_reg_4_ ( .D(n845), .CLK(Clk), .QN(n22) );
  fd1c2 register_register1_reg_3_ ( .D(n849), .CLK(Clk), .QN(n18) );
  fd1c2 register_register1_reg_2_ ( .D(n853), .CLK(Clk), .QN(n14) );
  fd1c2 register_register1_reg_1_ ( .D(n857), .CLK(Clk), .QN(n10) );
  fd1c2 register_register3_reg_0_ ( .D(n859), .CLK(Clk), .QN(n8) );
  fd1c2 register_register1_reg_0_ ( .D(n861), .CLK(Clk), .QN(n6) );
  fd1c2 register_register3_reg_30_ ( .D(n739), .CLK(Clk), .QN(n4) );
  fd1c2 register_register1_reg_30_ ( .D(n741), .CLK(Clk), .QN(n2) );
  fd1c2 register_register3_reg_31_ ( .D(n736), .CLK(Clk), .QN(n127) );
  fd1c2 register_register3_reg_27_ ( .D(n751), .CLK(Clk), .QN(n124) );
  fd1c2 register_register3_reg_28_ ( .D(n747), .CLK(Clk), .QN(n120) );
  fd1c2 register_register3_reg_29_ ( .D(n743), .CLK(Clk), .QN(n116) );
  fd1c2 register_register3_reg_26_ ( .D(n755), .CLK(Clk), .QN(n112) );
  fd1c2 register_register3_reg_25_ ( .D(n759), .CLK(Clk), .QN(n108) );
  fd1c2 register_register3_reg_24_ ( .D(n763), .CLK(Clk), .QN(n104) );
  fd1c2 register_register3_reg_23_ ( .D(n767), .CLK(Clk), .QN(n100) );
  fd1c2 register_register3_reg_22_ ( .D(n771), .CLK(Clk), .QN(n96) );
  fd1c2 register_register3_reg_21_ ( .D(n775), .CLK(Clk), .QN(n92) );
  fd1c2 register_register3_reg_20_ ( .D(n779), .CLK(Clk), .QN(n88) );
  fd1c2 register_register3_reg_19_ ( .D(n783), .CLK(Clk), .QN(n84) );
  fd1c2 register_register3_reg_18_ ( .D(n787), .CLK(Clk), .QN(n80) );
  fd1c2 register_register3_reg_17_ ( .D(n791), .CLK(Clk), .QN(n76) );
  fd1c2 register_register3_reg_16_ ( .D(n795), .CLK(Clk), .QN(n72) );
  fd1c2 register_register3_reg_15_ ( .D(n799), .CLK(Clk), .QN(n68) );
  fd1c2 register_register3_reg_14_ ( .D(n803), .CLK(Clk), .QN(n64) );
  fd1c2 register_register3_reg_13_ ( .D(n807), .CLK(Clk), .QN(n60) );
  fd1c2 register_register3_reg_12_ ( .D(n811), .CLK(Clk), .QN(n56) );
  fd1c2 register_register3_reg_11_ ( .D(n815), .CLK(Clk), .QN(n52) );
  fd1c2 register_register3_reg_10_ ( .D(n819), .CLK(Clk), .QN(n48) );
  fd1c2 register_register3_reg_9_ ( .D(n823), .CLK(Clk), .QN(n44) );
  fd1c2 register_register3_reg_8_ ( .D(n827), .CLK(Clk), .QN(n40) );
  fd1c2 register_register3_reg_7_ ( .D(n831), .CLK(Clk), .QN(n36) );
  fd1c2 register_register3_reg_6_ ( .D(n835), .CLK(Clk), .QN(n32) );
  fd1c2 register_register3_reg_5_ ( .D(n839), .CLK(Clk), .QN(n28) );
  fd1c2 register_register3_reg_4_ ( .D(n843), .CLK(Clk), .QN(n24) );
  fd1c2 register_register3_reg_3_ ( .D(n847), .CLK(Clk), .QN(n20) );
  fd1c2 register_register3_reg_2_ ( .D(n851), .CLK(Clk), .QN(n16) );
  fd1c2 register_register3_reg_1_ ( .D(n855), .CLK(Clk), .QN(n12) );
  fd1c2 register_register2_reg_31_ ( .D(n895), .CLK(Clk), .QN(n128) );
  fd1c2 register_register2_reg_27_ ( .D(n752), .CLK(Clk), .QN(n123) );
  fd1c2 register_register2_reg_28_ ( .D(n748), .CLK(Clk), .QN(n119) );
  fd1c2 register_register2_reg_29_ ( .D(n744), .CLK(Clk), .QN(n115) );
  fd1c2 register_register2_reg_26_ ( .D(n756), .CLK(Clk), .QN(n111) );
  fd1c2 register_register2_reg_25_ ( .D(n760), .CLK(Clk), .QN(n107) );
  fd1c2 register_register2_reg_24_ ( .D(n764), .CLK(Clk), .QN(n103) );
  fd1c2 register_register2_reg_23_ ( .D(n768), .CLK(Clk), .QN(n99) );
  fd1c2 register_register2_reg_22_ ( .D(n772), .CLK(Clk), .QN(n95) );
  fd1c2 register_register2_reg_21_ ( .D(n776), .CLK(Clk), .QN(n91) );
  fd1c2 register_register2_reg_20_ ( .D(n780), .CLK(Clk), .QN(n87) );
  fd1c2 register_register2_reg_19_ ( .D(n784), .CLK(Clk), .QN(n83) );
  fd1c2 register_register2_reg_18_ ( .D(n788), .CLK(Clk), .QN(n79) );
  fd1c2 register_register2_reg_17_ ( .D(n792), .CLK(Clk), .QN(n75) );
  fd1c2 register_register2_reg_16_ ( .D(n796), .CLK(Clk), .QN(n71) );
  fd1c2 register_register2_reg_15_ ( .D(n800), .CLK(Clk), .QN(n67) );
  fd1c2 register_register2_reg_14_ ( .D(n804), .CLK(Clk), .QN(n63) );
  fd1c2 register_register2_reg_13_ ( .D(n808), .CLK(Clk), .QN(n59) );
  fd1c2 register_register2_reg_12_ ( .D(n812), .CLK(Clk), .QN(n55) );
  fd1c2 register_register2_reg_11_ ( .D(n816), .CLK(Clk), .QN(n51) );
  fd1c2 register_register2_reg_9_ ( .D(n824), .CLK(Clk), .QN(n43) );
  fd1c2 register_register2_reg_8_ ( .D(n828), .CLK(Clk), .QN(n39) );
  fd1c2 register_register2_reg_7_ ( .D(n832), .CLK(Clk), .QN(n35) );
  fd1c2 register_register2_reg_6_ ( .D(n836), .CLK(Clk), .QN(n31) );
  fd1c2 register_register2_reg_4_ ( .D(n844), .CLK(Clk), .QN(n23) );
  fd1c2 register_register2_reg_3_ ( .D(n848), .CLK(Clk), .QN(n19) );
  fd1c2 register_register2_reg_2_ ( .D(n852), .CLK(Clk), .QN(n15) );
  fd1c2 register_register2_reg_1_ ( .D(n856), .CLK(Clk), .QN(n11) );
  fd1c2 register_register2_reg_0_ ( .D(n860), .CLK(Clk), .QN(n7) );
  fd1c2 register_register2_reg_30_ ( .D(n740), .CLK(Clk), .QN(n3) );
  fd1c2 register_register0_reg_31_ ( .D(n738), .CLK(Clk), .QN(n125) );
  fd1c2 register_register0_reg_27_ ( .D(n754), .CLK(Clk), .QN(n121) );
  fd1c2 register_register0_reg_28_ ( .D(n750), .CLK(Clk), .QN(n117) );
  fd1c2 register_register0_reg_29_ ( .D(n746), .CLK(Clk), .QN(n113) );
  fd1c2 register_register0_reg_26_ ( .D(n758), .CLK(Clk), .QN(n109) );
  fd1c2 register_register0_reg_25_ ( .D(n762), .CLK(Clk), .QN(n105) );
  fd1c2 register_register0_reg_24_ ( .D(n766), .CLK(Clk), .QN(n101) );
  fd1c2 register_register0_reg_23_ ( .D(n770), .CLK(Clk), .QN(n97) );
  fd1c2 register_register0_reg_22_ ( .D(n774), .CLK(Clk), .QN(n93) );
  fd1c2 register_register0_reg_21_ ( .D(n778), .CLK(Clk), .QN(n89) );
  fd1c2 register_register0_reg_20_ ( .D(n782), .CLK(Clk), .QN(n85) );
  fd1c2 register_register0_reg_19_ ( .D(n786), .CLK(Clk), .QN(n81) );
  fd1c2 register_register0_reg_18_ ( .D(n790), .CLK(Clk), .QN(n77) );
  fd1c2 register_register0_reg_17_ ( .D(n794), .CLK(Clk), .QN(n73) );
  fd1c2 register_register0_reg_16_ ( .D(n798), .CLK(Clk), .QN(n69) );
  fd1c2 register_register0_reg_15_ ( .D(n802), .CLK(Clk), .QN(n65) );
  fd1c2 register_register0_reg_14_ ( .D(n806), .CLK(Clk), .QN(n61) );
  fd1c2 register_register0_reg_13_ ( .D(n810), .CLK(Clk), .QN(n57) );
  fd1c2 register_register0_reg_12_ ( .D(n814), .CLK(Clk), .QN(n53) );
  fd1c2 register_register0_reg_11_ ( .D(n818), .CLK(Clk), .QN(n49) );
  fd1c2 register_register2_reg_10_ ( .D(n820), .CLK(Clk), .QN(n47) );
  fd1c2 register_register0_reg_10_ ( .D(n822), .CLK(Clk), .QN(n45) );
  fd1c2 register_register0_reg_9_ ( .D(n826), .CLK(Clk), .QN(n41) );
  fd1c2 register_register0_reg_8_ ( .D(n830), .CLK(Clk), .QN(n37) );
  fd1c2 register_register0_reg_7_ ( .D(n834), .CLK(Clk), .QN(n33) );
  fd1c2 register_register0_reg_6_ ( .D(n838), .CLK(Clk), .QN(n29) );
  fd1c2 register_register2_reg_5_ ( .D(n840), .CLK(Clk), .QN(n27) );
  fd1c2 register_register0_reg_5_ ( .D(n842), .CLK(Clk), .QN(n25) );
  fd1c2 register_register0_reg_4_ ( .D(n846), .CLK(Clk), .QN(n21) );
  fd1c2 register_register0_reg_3_ ( .D(n850), .CLK(Clk), .QN(n17) );
  fd1c2 register_register0_reg_2_ ( .D(n854), .CLK(Clk), .QN(n13) );
  fd1c2 register_register0_reg_1_ ( .D(n858), .CLK(Clk), .QN(n9) );
  fd1c2 register_register0_reg_0_ ( .D(n862), .CLK(Clk), .QN(n5) );
  fd1c2 register_register0_reg_30_ ( .D(n742), .CLK(Clk), .QN(n1) );
  fd1a2 cntrl_ALUSelB_reg_0_ ( .D(cntrl_N109), .CLK(Clk), .Q(ALUSelB[0]) );
  fd1a2 cntrl_ALUOp_reg_0_ ( .D(cntrl_N111), .CLK(Clk), .Q(ALUOp[0]) );
  fd1a2 cntrl_MemtoReg_reg ( .D(n155), .CLK(Clk), .Q(MemToReg) );
  fd1a2 cntrl_state_reg_9_ ( .D(cntrl_N106), .CLK(Clk), .Q(cntrl_state_9_) );
  fd1a2 cntrl_PCSource_reg_0_ ( .D(cntrl_N111), .CLK(Clk), .Q(PCSource[0]) );
  fd1a2 cntrl_state_reg_10_ ( .D(n900), .CLK(Clk), .Q(cntrl_state_10_) );
  fde1a2 Instruction_reg_30_ ( .D(MemData[30]), .E(n978), .CLK(Clk), .Q(
        Instruction_30) );
  fde1a2 Instruction_reg_3_ ( .D(MemData[3]), .E(n978), .CLK(Clk), .Q(
        Instruction[3]) );
  fde1a2 Instruction_reg_4_ ( .D(MemData[4]), .E(n977), .CLK(Clk), .Q(
        Instruction[4]) );
  fde1a2 Instruction_reg_6_ ( .D(MemData[6]), .E(n977), .CLK(Clk), .Q(
        Instruction[6]) );
  fde1a2 Instruction_reg_7_ ( .D(MemData[7]), .E(n977), .CLK(Clk), .Q(
        Instruction[7]) );
  fde1a2 Instruction_reg_8_ ( .D(MemData[8]), .E(n977), .CLK(Clk), .Q(
        Instruction[8]) );
  fde1a2 Instruction_reg_9_ ( .D(MemData[9]), .E(n977), .CLK(Clk), .Q(
        Instruction[9]) );
  fde1a2 Instruction_reg_13_ ( .D(MemData[13]), .E(n977), .CLK(Clk), .Q(
        Instruction[13]) );
  fde1a2 Instruction_reg_14_ ( .D(MemData[14]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction[14]) );
  fdm5a2 cntrl_PCSource_reg_1_ ( .D0(n142), .D1(n972), .D2(n144), .S0(
        cntrl_state_10_), .S1(n900), .CLK(Clk), .Q(PCSource[1]) );
  fde1a2 Instruction_reg_28_ ( .D(MemData[28]), .E(n978), .CLK(Clk), .Q(
        Instruction_28) );
  fde1a2 Instruction_reg_10_ ( .D(MemData[10]), .E(n977), .CLK(Clk), .Q(
        Instruction[10]) );
  fde1a2 Instruction_reg_31_ ( .D(MemData[31]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction_31) );
  fde1a2 Instruction_reg_26_ ( .D(MemData[26]), .E(n978), .CLK(Clk), .Q(
        Instruction_26) );
  fd1a2 cntrl_RegDst_reg ( .D(cntrl_N114), .CLK(Clk), .Q(RegDst) );
  fde1a2 Instruction_reg_15_ ( .D(MemData[15]), .E(n978), .CLK(Clk), .Q(
        Instruction[15]) );
  fdm5a2 cntrl_state_reg_8_ ( .D0(n142), .D1(cntrl_state_1_), .D2(n142), .S0(
        n145), .S1(Reset), .CLK(Clk), .Q(cntrl_state_8_) );
  fdm5a2 cntrl_RegWrite_reg ( .D0(n142), .D1(n419), .D2(n144), .S0(n155), .S1(
        n156), .CLK(Clk), .Q(RegWrite) );
  fdm5a2 cntrl_state_reg_3_ ( .D0(n142), .D1(cntrl_state_2_), .D2(n142), .S0(
        n971), .S1(n140), .CLK(Clk), .Q(cntrl_state_3_) );
  fd1a2 cntrl_state_reg_6_ ( .D(n896), .CLK(Clk), .Q(cntrl_state_6_) );
  fdm5a2 cntrl_state_reg_0_ ( .D0(cntrl_state_7_), .D1(n144), .D2(n144), .S0(
        n426), .S1(Reset), .CLK(Clk), .Q(cntrl_state_0_) );
  fde1a2 Instruction_reg_1_ ( .D(MemData[1]), .E(n978), .CLK(Clk), .Q(
        Instruction[1]) );
  fde1a2 Instruction_reg_29_ ( .D(MemData[29]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction_29) );
  fde1a2 Instruction_reg_11_ ( .D(MemData[11]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction[11]) );
  fde1a2 Instruction_reg_12_ ( .D(MemData[12]), .E(n978), .CLK(Clk), .Q(
        Instruction[12]) );
  fde1a2 Instruction_reg_2_ ( .D(MemData[2]), .E(n978), .CLK(Clk), .Q(
        Instruction[2]) );
  fd2a2 PC_reg_27_ ( .D(n867), .CLK(Clk), .CLR(n972), .Q(PC[27]) );
  fd2a2 PC_reg_26_ ( .D(n868), .CLK(Clk), .CLR(n972), .Q(PC[26]) );
  fd2a2 PC_reg_25_ ( .D(n869), .CLK(Clk), .CLR(n972), .Q(PC[25]) );
  fd2a2 PC_reg_24_ ( .D(n870), .CLK(Clk), .CLR(n972), .Q(PC[24]) );
  fd2a2 PC_reg_23_ ( .D(n871), .CLK(Clk), .CLR(n972), .Q(PC[23]) );
  fd2a2 PC_reg_22_ ( .D(n872), .CLK(Clk), .CLR(n972), .Q(PC[22]) );
  fd2a2 PC_reg_21_ ( .D(n873), .CLK(Clk), .CLR(n972), .Q(PC[21]) );
  fd2a2 PC_reg_20_ ( .D(n874), .CLK(Clk), .CLR(n157), .Q(PC[20]) );
  fd2a2 PC_reg_19_ ( .D(n875), .CLK(Clk), .CLR(n157), .Q(PC[19]) );
  fd2a2 PC_reg_18_ ( .D(n876), .CLK(Clk), .CLR(n157), .Q(PC[18]) );
  fd2a2 PC_reg_17_ ( .D(n877), .CLK(Clk), .CLR(n971), .Q(PC[17]) );
  fd2a2 PC_reg_16_ ( .D(n878), .CLK(Clk), .CLR(n972), .Q(PC[16]) );
  fd2a2 PC_reg_15_ ( .D(n879), .CLK(Clk), .CLR(n971), .Q(PC[15]) );
  fd2a2 PC_reg_14_ ( .D(n880), .CLK(Clk), .CLR(n972), .Q(PC[14]) );
  fd2a2 PC_reg_13_ ( .D(n881), .CLK(Clk), .CLR(n971), .Q(PC[13]) );
  fd2a2 PC_reg_12_ ( .D(n882), .CLK(Clk), .CLR(n972), .Q(PC[12]) );
  fd2a2 PC_reg_11_ ( .D(n883), .CLK(Clk), .CLR(n971), .Q(PC[11]) );
  fd2a2 PC_reg_10_ ( .D(n884), .CLK(Clk), .CLR(n971), .Q(PC[10]) );
  fd2a2 PC_reg_9_ ( .D(n885), .CLK(Clk), .CLR(n971), .Q(PC[9]) );
  fd2a2 PC_reg_8_ ( .D(n886), .CLK(Clk), .CLR(n972), .Q(PC[8]) );
  fd2a2 PC_reg_7_ ( .D(n887), .CLK(Clk), .CLR(n972), .Q(PC[7]) );
  fd2a2 PC_reg_6_ ( .D(n888), .CLK(Clk), .CLR(n972), .Q(PC[6]) );
  fd2a2 PC_reg_5_ ( .D(n889), .CLK(Clk), .CLR(n971), .Q(PC[5]) );
  fd2a2 PC_reg_4_ ( .D(n890), .CLK(Clk), .CLR(n157), .Q(PC[4]) );
  fd2a2 PC_reg_3_ ( .D(n891), .CLK(Clk), .CLR(n972), .Q(PC[3]) );
  fd2a2 PC_reg_1_ ( .D(n893), .CLK(Clk), .CLR(n972), .Q(PC[1]) );
  fd2a2 PC_reg_2_ ( .D(n892), .CLK(Clk), .CLR(n971), .Q(PC[2]) );
  fd2a2 PC_reg_0_ ( .D(n894), .CLK(Clk), .CLR(n971), .Q(PC[0]) );
  fde1a2 Instruction_reg_0_ ( .D(MemData[0]), .E(n978), .CLK(Clk), .Q(
        Instruction[0]) );
  fde1a2 Instruction_reg_27_ ( .D(MemData[27]), .E(IRWrite), .CLK(Clk), .Q(
        Instruction_27) );
  fde1a2 Instruction_reg_22_ ( .D(MemData[22]), .E(IRWrite), .CLK(Clk), .Q(
        Read1RegSel[1]) );
  fd1a2 cntrl_ALUOp_reg_1_ ( .D(n156), .CLK(Clk), .Q(ALUOp[1]) );
  fd2a2 PC_reg_31_ ( .D(n863), .CLK(Clk), .CLR(n157), .Q(PC[31]) );
  fd2a2 PC_reg_30_ ( .D(n864), .CLK(Clk), .CLR(n972), .Q(PC[30]) );
  fd2a2 PC_reg_29_ ( .D(n865), .CLK(Clk), .CLR(n971), .Q(PC[29]) );
  fd2a2 PC_reg_28_ ( .D(n866), .CLK(Clk), .CLR(n157), .Q(PC[28]) );
  fde1a2 Instruction_reg_16_ ( .D(MemData[16]), .E(n977), .CLK(Clk), .Q(
        Read2RegSel[0]) );
  fde1a2 Instruction_reg_17_ ( .D(MemData[17]), .E(IRWrite), .CLK(Clk), .Q(
        Read2RegSel[1]) );
  fd1a2 cntrl_state_reg_1_ ( .D(n899), .CLK(Clk), .Q(cntrl_state_1_) );
  fde1a2 Instruction_reg_5_ ( .D(MemData[5]), .E(n977), .CLK(Clk), .Q(
        Instruction[5]) );
  fde1a2 Instruction_reg_21_ ( .D(MemData[21]), .E(IRWrite), .CLK(Clk), .Q(
        Read1RegSel[0]) );
  fd1a2 cntrl_state_reg_7_ ( .D(n156), .CLK(Clk), .Q(cntrl_state_7_) );
  fd1a2 cntrl_state_reg_2_ ( .D(n898), .CLK(Clk), .Q(cntrl_state_2_) );
  fdm5a2 cntrl_ALUSelB_reg_1_ ( .D0(cntrl_state_2_), .D1(n144), .D2(n142), 
        .S0(cntrl_state_1_), .S1(Reset), .CLK(Clk), .Q(ALUSelB[1]) );
  xor2a2 DP_OP_100J1_124_3689_U65 ( .A(alu_MuxB_1_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n66) );
  xor2a2 DP_OP_100J1_124_3689_U64 ( .A(alu_MuxB_2_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n65) );
  xor2a2 DP_OP_100J1_124_3689_U63 ( .A(alu_MuxB_3_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n64) );
  xor2a2 DP_OP_100J1_124_3689_U62 ( .A(alu_MuxB_4_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n63) );
  xor2a2 DP_OP_100J1_124_3689_U61 ( .A(alu_MuxB_5_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n62) );
  xor2a2 DP_OP_100J1_124_3689_U60 ( .A(alu_MuxB_6_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n61) );
  xor2a2 DP_OP_100J1_124_3689_U59 ( .A(alu_MuxB_7_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n60) );
  xor2a2 DP_OP_100J1_124_3689_U58 ( .A(alu_MuxB_8_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n59) );
  xor2a2 DP_OP_100J1_124_3689_U57 ( .A(alu_MuxB_9_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n58) );
  xor2a2 DP_OP_100J1_124_3689_U56 ( .A(alu_MuxB_10_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n57) );
  xor2a2 DP_OP_100J1_124_3689_U55 ( .A(alu_MuxB_11_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n56) );
  xor2a2 DP_OP_100J1_124_3689_U54 ( .A(alu_MuxB_12_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n55) );
  xor2a2 DP_OP_100J1_124_3689_U53 ( .A(alu_MuxB_13_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n54) );
  xor2a2 DP_OP_100J1_124_3689_U52 ( .A(alu_MuxB_14_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n53) );
  xor2a2 DP_OP_100J1_124_3689_U51 ( .A(alu_MuxB_15_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n52) );
  xor2a2 DP_OP_100J1_124_3689_U35 ( .A(alu_MuxB_31_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n36) );
  xor2a2 DP_OP_100J1_124_3689_U36 ( .A(alu_MuxB_30_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n37) );
  xor2a2 DP_OP_100J1_124_3689_U37 ( .A(alu_MuxB_29_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n38) );
  xor2a2 DP_OP_100J1_124_3689_U38 ( .A(alu_MuxB_28_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n39) );
  xor2a2 DP_OP_100J1_124_3689_U39 ( .A(alu_MuxB_27_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n40) );
  xor2a2 DP_OP_100J1_124_3689_U40 ( .A(alu_MuxB_26_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n41) );
  xor2a2 DP_OP_100J1_124_3689_U41 ( .A(alu_MuxB_25_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n42) );
  xor2a2 DP_OP_100J1_124_3689_U42 ( .A(alu_MuxB_24_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n43) );
  xor2a2 DP_OP_100J1_124_3689_U43 ( .A(alu_MuxB_23_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n44) );
  xor2a2 DP_OP_100J1_124_3689_U44 ( .A(alu_MuxB_22_), .B(n927), .Y(
        DP_OP_100J1_124_3689_n45) );
  xor2a2 DP_OP_100J1_124_3689_U45 ( .A(alu_MuxB_21_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n46) );
  xor2a2 DP_OP_100J1_124_3689_U46 ( .A(alu_MuxB_20_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n47) );
  xor2a2 DP_OP_100J1_124_3689_U47 ( .A(alu_MuxB_19_), .B(n926), .Y(
        DP_OP_100J1_124_3689_n48) );
  xor2a2 DP_OP_100J1_124_3689_U48 ( .A(alu_MuxB_18_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n49) );
  xor2a2 DP_OP_100J1_124_3689_U49 ( .A(alu_MuxB_17_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n50) );
  xor2a2 DP_OP_100J1_124_3689_U50 ( .A(alu_MuxB_16_), .B(
        DP_OP_100J1_124_3689_n100), .Y(DP_OP_100J1_124_3689_n51) );
  mx2d0 U1073 ( .D0(Read2RegSel[0]), .D1(Instruction[11]), .S(RegDst), .Y(
        n1441) );
  inv1a1 U1074 ( .A(Read2RegSel[1]), .Y(n1151) );
  inv1a1 U1075 ( .A(Read2RegSel[0]), .Y(n1150) );
  mx2d0 U1076 ( .D0(Read2RegSel[1]), .D1(Instruction[12]), .S(RegDst), .Y(
        n1442) );
  and2c0 U1077 ( .A(Instruction[2]), .B(n1022), .Y(n1018) );
  or2c0 U1078 ( .A(ALUOp[1]), .B(Instruction[1]), .Y(n1159) );
  inv1a1 U1079 ( .A(Instruction[5]), .Y(n1022) );
  or2c0 U1080 ( .A(ALUOp[1]), .B(n1148), .Y(n1170) );
  inv1a1 U1081 ( .A(Instruction[2]), .Y(n1149) );
  inv1a1 U1082 ( .A(Instruction[1]), .Y(n1148) );
  nor2a0 U1083 ( .A(n1159), .B(n1149), .Y(n1298) );
  inv1a1 U1084 ( .A(n1298), .Y(n1345) );
  ao1f1 U1085 ( .A(n1330), .B(n87), .C(n1225), .Y(WriteData[20]) );
  ao1f1 U1086 ( .A(n1330), .B(n91), .C(n1237), .Y(WriteData[21]) );
  ao1f1 U1087 ( .A(n1330), .B(n99), .C(n1249), .Y(WriteData[23]) );
  oa1d1 U1088 ( .A(cntrl_state_6_), .B(cntrl_state_7_), .C(Reset), .Y(
        cntrl_N114) );
  and2c0 U1089 ( .A(Reset), .B(n1354), .Y(n155) );
  and2b1 U1090 ( .B(Instruction_27), .A(n1359), .Y(n900) );
  or2c0 U1091 ( .A(n1441), .B(RegWrite), .Y(n1440) );
  ao7g0 U1092 ( .A(n935), .B(n121), .C(n933), .D(n122), .E(n937), .F(n124), 
        .Y(n903) );
  ao1c0 U1093 ( .A(n1330), .B(n123), .C(n903), .Y(WriteData[27]) );
  ao7g0 U1094 ( .A(n935), .B(n117), .C(n933), .D(n118), .E(n937), .F(n120), 
        .Y(n904) );
  ao1c0 U1095 ( .A(n1330), .B(n119), .C(n904), .Y(WriteData[28]) );
  nand3b0 U1096 ( .A(n973), .B(Read1RegSel[0]), .C(Read1RegSel[1]), .Y(n1339)
         );
  ao4d0 U1097 ( .B(ALUSelB[1]), .A(Instruction[0]), .D(n929), .C(WriteData[0]), 
        .Y(n921) );
  ao7g0 U1098 ( .A(n935), .B(n113), .C(n933), .D(n114), .E(n937), .F(n116), 
        .Y(n905) );
  ao1c0 U1099 ( .A(n939), .B(n115), .C(n905), .Y(WriteData[29]) );
  nand2b1 U1100 ( .A(Read1RegSel[0]), .B(n1154), .Y(n1011) );
  and2b1 U1101 ( .B(WriteData[5]), .A(n930), .Y(n1126) );
  ao7g0 U1102 ( .A(n934), .B(n1), .C(n932), .D(n2), .E(n936), .F(n4), .Y(n906)
         );
  ao1c0 U1103 ( .A(n1330), .B(n3), .C(n906), .Y(WriteData[30]) );
  nand2a0 U1104 ( .A(n1354), .B(n1355), .Y(n907) );
  or6a1 U1105 ( .A(n907), .B(n426), .C(cntrl_state_6_), .D(cntrl_state_7_), 
        .E(cntrl_state_8_), .F(cntrl_state_3_), .Y(n908) );
  ao4e0 U1106 ( .B(cntrl_state_0_), .A(Reset), .C(n1356), .D(n908), .Y(n899)
         );
  inv1a0 U1107 ( .A(n957), .Y(n909) );
  oa7g0 U1108 ( .A(n909), .B(Instruction[0]), .C(n1437), .D(PC[0]), .E(
        TargetReg[0]), .F(n959), .Y(n910) );
  ao1d1 U1109 ( .A(WriteAdd[0]), .B(n960), .C(n910), .Y(n894) );
  mx2d0 U1110 ( .D0(n926), .D1(alu_MuxA_0_), .S(n924), .Y(
        DP_OP_100J1_124_3689_n31) );
  inv1a0 U1111 ( .A(alu_MuxA_0_), .Y(n911) );
  mx2d0 U1112 ( .D0(n911), .D1(alu_MuxA_0_), .S(n924), .Y(C55_DATA6_0) );
  ao7g0 U1113 ( .A(n934), .B(n125), .C(n932), .D(n126), .E(n937), .F(n127), 
        .Y(n912) );
  ao1c0 U1114 ( .A(n1330), .B(n128), .C(n912), .Y(WriteData[31]) );
  and2c0 U1115 ( .A(Instruction_27), .B(Instruction_29), .Y(n913) );
  nand3a1 U1116 ( .A(n913), .B(n1351), .C(Instruction_28), .Y(n914) );
  and2c0 U1117 ( .A(Instruction_30), .B(n914), .Y(n145) );
  oa4f0 U1118 ( .A(n1143), .B(alu_MuxB_4_), .C(n1132), .D(alu_MuxB_6_), .Y(
        n915) );
  ao1f1 U1119 ( .A(alu_MuxA_5_), .B(n953), .C(n948), .Y(n916) );
  oa4f0 U1120 ( .A(n931), .B(C55_DATA6_5), .C(alu_MuxB_5_), .D(n916), .Y(n917)
         );
  nand2a0 U1121 ( .A(alu_MuxB_5_), .B(n947), .Y(n918) );
  ao2i0 U1122 ( .A(n955), .B(alu_MuxB_5_), .C(n949), .D(n918), .Y(n919) );
  nand2a0 U1123 ( .A(alu_MuxA_5_), .B(n919), .Y(n920) );
  nand3a1 U1124 ( .A(n920), .B(n915), .C(n917), .Y(WriteAdd[5]) );
  buf1a2 U1125 ( .A(n1438), .Y(n959) );
  or2c0 U1126 ( .A(MemToReg), .B(n157), .Y(n922) );
  inv1a1 U1127 ( .A(n1013), .Y(n930) );
  buf1a2 U1128 ( .A(n1479), .Y(n968) );
  buf1a2 U1129 ( .A(n1480), .Y(n970) );
  inv1a1 U1130 ( .A(n1434), .Y(n957) );
  buf1a2 U1131 ( .A(n1330), .Y(n939) );
  nand2a1 U1132 ( .A(Read2RegSel[0]), .B(Read2RegSel[1]), .Y(n1328) );
  ao1a2 U1133 ( .A(Instruction[5]), .B(ALUSelB[1]), .C(n1126), .Y(alu_MuxB_5_)
         );
  inv1a4 U1134 ( .A(n922), .Y(n923) );
  inv1a1 U1135 ( .A(n921), .Y(n924) );
  oa4f1 U1136 ( .A(MemData[29]), .B(n962), .C(n1475), .D(WriteAdd[29]), .Y(
        n1474) );
  ao2i1 U1137 ( .A(n1116), .B(n1146), .C(n1103), .D(n1102), .Y(WriteAdd[29])
         );
  oa4f1 U1138 ( .A(MemData[27]), .B(n962), .C(n1475), .D(WriteAdd[27]), .Y(
        n1472) );
  ao2i1 U1139 ( .A(n1096), .B(n1146), .C(n1095), .D(n1094), .Y(WriteAdd[27])
         );
  oa4f1 U1140 ( .A(MemData[26]), .B(n962), .C(n1475), .D(WriteAdd[26]), .Y(
        n1471) );
  ao2i1 U1141 ( .A(n1092), .B(n1146), .C(n1091), .D(n1090), .Y(WriteAdd[26])
         );
  oa4f1 U1142 ( .A(MemData[23]), .B(n962), .C(n1475), .D(WriteAdd[23]), .Y(
        n1468) );
  ao2i1 U1143 ( .A(n1080), .B(n1146), .C(n1079), .D(n1078), .Y(WriteAdd[23])
         );
  oa4f1 U1144 ( .A(MemData[21]), .B(n962), .C(n961), .D(WriteAdd[21]), .Y(
        n1466) );
  ao2i1 U1145 ( .A(n1072), .B(n1146), .C(n1071), .D(n1070), .Y(WriteAdd[21])
         );
  oa4f1 U1146 ( .A(MemData[20]), .B(n923), .C(n961), .D(WriteAdd[20]), .Y(
        n1465) );
  and3d1 U1147 ( .A(WriteAdd[20]), .B(WriteAdd[19]), .C(n1364), .Y(n1374) );
  ao2i1 U1148 ( .A(n1068), .B(n1146), .C(n1067), .D(n1066), .Y(WriteAdd[20])
         );
  oa4f1 U1149 ( .A(MemData[19]), .B(n962), .C(n961), .D(WriteAdd[19]), .Y(
        n1464) );
  ao2i1 U1150 ( .A(n1061), .B(n1146), .C(n1060), .D(n1059), .Y(WriteAdd[19])
         );
  oa4f1 U1151 ( .A(MemData[17]), .B(n962), .C(n961), .D(WriteAdd[17]), .Y(
        n1462) );
  ao2i1 U1152 ( .A(n1053), .B(n1146), .C(n1052), .D(n1051), .Y(WriteAdd[17])
         );
  ao2i1 U1153 ( .A(n1116), .B(n1135), .C(n1115), .D(n1114), .Y(WriteAdd[31])
         );
  oa4f1 U1154 ( .A(MemData[31]), .B(n923), .C(n1475), .D(WriteAdd[31]), .Y(
        n1481) );
  oa4f1 U1155 ( .A(MemData[7]), .B(n962), .C(n961), .D(WriteAdd[7]), .Y(n1452)
         );
  ao2i1 U1156 ( .A(n1136), .B(n1135), .C(n1134), .D(n1133), .Y(WriteAdd[7]) );
  oa4f1 U1157 ( .A(MemData[6]), .B(n923), .C(n1475), .D(WriteAdd[6]), .Y(n1451) );
  and3d1 U1158 ( .A(WriteAdd[6]), .B(WriteAdd[5]), .C(n1371), .Y(n1372) );
  or4e1 U1159 ( .A(n1130), .B(n1129), .C(n1128), .D(n1127), .Y(WriteAdd[6]) );
  oa4f1 U1160 ( .A(MemData[5]), .B(n923), .C(n1475), .D(WriteAdd[5]), .Y(n1450) );
  oa4f1 U1161 ( .A(MemData[1]), .B(n923), .C(n961), .D(WriteAdd[1]), .Y(n1446)
         );
  ao2i1 U1162 ( .A(n1135), .B(n921), .C(n1064), .D(n1063), .Y(WriteAdd[1]) );
  ao2i1 U1163 ( .A(n1111), .B(n1146), .C(n1110), .D(n1109), .Y(WriteAdd[30])
         );
  oa4f1 U1164 ( .A(MemData[30]), .B(n962), .C(n961), .D(WriteAdd[30]), .Y(
        n1477) );
  oa4f1 U1165 ( .A(MemData[18]), .B(n923), .C(n1475), .D(WriteAdd[18]), .Y(
        n1463) );
  ao2i1 U1166 ( .A(n1057), .B(n1146), .C(n1056), .D(n1055), .Y(WriteAdd[18])
         );
  oa4f1 U1167 ( .A(MemData[2]), .B(n962), .C(n961), .D(WriteAdd[2]), .Y(n1447)
         );
  ao2i1 U1168 ( .A(n1107), .B(n1135), .C(n1106), .D(n1105), .Y(WriteAdd[2]) );
  ao2i1 U1169 ( .A(n1088), .B(n1146), .C(n1087), .D(n1086), .Y(WriteAdd[25])
         );
  nor2a0 U1170 ( .A(WriteAdd[26]), .B(WriteAdd[25]), .Y(n1361) );
  ao2i1 U1171 ( .A(n1045), .B(n1146), .C(n1044), .D(n1043), .Y(WriteAdd[15])
         );
  ao2i1 U1172 ( .A(n1041), .B(n1146), .C(n1040), .D(n1039), .Y(WriteAdd[14])
         );
  and3d1 U1173 ( .A(WriteAdd[14]), .B(WriteAdd[13]), .C(n1367), .Y(n1373) );
  ao2i1 U1174 ( .A(n1037), .B(n1135), .C(n1036), .D(n1035), .Y(WriteAdd[13])
         );
  ao2i1 U1175 ( .A(n1147), .B(n1146), .C(n1145), .D(n1144), .Y(WriteAdd[9]) );
  ao2i1 U1176 ( .A(n1120), .B(n1135), .C(n1119), .D(n1118), .Y(WriteAdd[3]) );
  ao2i1 U1177 ( .A(n1033), .B(n1135), .C(n1032), .D(n1031), .Y(WriteAdd[12])
         );
  ao2i1 U1178 ( .A(n1100), .B(n1146), .C(n1099), .D(n1098), .Y(WriteAdd[28])
         );
  ao2i1 U1179 ( .A(n1084), .B(n1146), .C(n1083), .D(n1082), .Y(WriteAdd[24])
         );
  ao2i1 U1180 ( .A(n1049), .B(n1146), .C(n1048), .D(n1047), .Y(WriteAdd[16])
         );
  ao2i1 U1181 ( .A(n1140), .B(n1146), .C(n1139), .D(n1138), .Y(WriteAdd[8]) );
  ao2i1 U1182 ( .A(n1107), .B(n1146), .C(n1021), .D(n1020), .Y(WriteAdd[0]) );
  ao4f1 U1183 ( .A(n1014), .B(n930), .C(n1015), .D(n1149), .Y(alu_MuxB_2_) );
  oa1d2 U1184 ( .A(n1377), .B(n1376), .C(PCWrite), .Y(n1437) );
  inv1a1 U1185 ( .A(Reset), .Y(n157) );
  inv1a1 U1186 ( .A(n957), .Y(n956) );
  ao4f1 U1187 ( .A(n1016), .B(n930), .C(n1015), .D(n1148), .Y(alu_MuxB_1_) );
  oa4f1 U1188 ( .A(MemData[10]), .B(n962), .C(n961), .D(WriteAdd[10]), .Y(
        n1455) );
  nand3a1 U1189 ( .A(n1026), .B(n1025), .C(n1024), .Y(WriteAdd[10]) );
  oa4f1 U1190 ( .A(MemData[4]), .B(n962), .C(n1475), .D(WriteAdd[4]), .Y(n1449) );
  or4e1 U1191 ( .A(n1125), .B(n1124), .C(n1123), .D(n1122), .Y(WriteAdd[4]) );
  ao2i1 U1192 ( .A(n1076), .B(n1146), .C(n1075), .D(n1074), .Y(WriteAdd[22])
         );
  ao2i1 U1193 ( .A(n1147), .B(n1135), .C(n1029), .D(n1028), .Y(WriteAdd[11])
         );
  buf1a2 U1194 ( .A(n1012), .Y(n925) );
  nand2a1 U1195 ( .A(ALUSelB[1]), .B(Instruction[15]), .Y(n1012) );
  buf1a2 U1196 ( .A(n1476), .Y(n963) );
  buf1a2 U1197 ( .A(n1478), .Y(n965) );
  ao1a2 U1198 ( .A(n1018), .B(n1017), .C(ALUOp[0]), .Y(
        DP_OP_100J1_124_3689_n100) );
  buf1a4 U1199 ( .A(n1344), .Y(n949) );
  or2c0 U1200 ( .A(Instruction[0]), .B(ALUOp[1]), .Y(n1344) );
  inv1a0 U1201 ( .A(n419), .Y(n140) );
  and2c0 U1202 ( .A(n1358), .B(n1357), .Y(n898) );
  oa3h1 U1203 ( .A(n1442), .B(RegWrite), .C(n1443), .D(Reset), .Y(n1479) );
  and2c0 U1204 ( .A(Reset), .B(n1353), .Y(cntrl_N116) );
  nand2a0 U1205 ( .A(n1348), .B(n157), .Y(cntrl_N104) );
  and2a2 U1206 ( .A(cntrl_state_3_), .B(n972), .Y(n897) );
  oa3h1 U1207 ( .A(RegWrite), .B(n1444), .C(n1443), .D(Reset), .Y(n1480) );
  inv1a0 U1208 ( .A(n1441), .Y(n1443) );
  nand2a0 U1209 ( .A(n1389), .B(n1388), .Y(n888) );
  nand2a0 U1210 ( .A(n1391), .B(n1390), .Y(n887) );
  nand2a0 U1211 ( .A(n1385), .B(n1384), .Y(n890) );
  nand2a0 U1212 ( .A(n1393), .B(n1392), .Y(n886) );
  nand2a0 U1213 ( .A(n1395), .B(n1394), .Y(n885) );
  nand2a0 U1214 ( .A(n1383), .B(n1382), .Y(n891) );
  nand2a0 U1215 ( .A(n1397), .B(n1396), .Y(n884) );
  nand2a0 U1216 ( .A(n1399), .B(n1398), .Y(n883) );
  nand2a0 U1217 ( .A(n1439), .B(WriteAdd[1]), .Y(n1378) );
  nand2a0 U1218 ( .A(n1401), .B(n1400), .Y(n882) );
  nand2a0 U1219 ( .A(n1403), .B(n1402), .Y(n881) );
  nand2a0 U1220 ( .A(n1405), .B(n1404), .Y(n880) );
  nand2a0 U1221 ( .A(n1407), .B(n1406), .Y(n879) );
  nand2a0 U1222 ( .A(n1409), .B(n1408), .Y(n878) );
  nand2a0 U1223 ( .A(n1411), .B(n1410), .Y(n877) );
  nand2a0 U1224 ( .A(n1413), .B(n1412), .Y(n876) );
  nand2a0 U1225 ( .A(n1415), .B(n1414), .Y(n875) );
  and2a2 U1226 ( .A(cntrl_state_6_), .B(n971), .Y(n156) );
  nand2a0 U1227 ( .A(n1417), .B(n1416), .Y(n874) );
  nand2a0 U1228 ( .A(n1419), .B(n1418), .Y(n873) );
  nand2a0 U1229 ( .A(n1421), .B(n1420), .Y(n872) );
  nand2a0 U1230 ( .A(n1423), .B(n1422), .Y(n871) );
  nand2a0 U1231 ( .A(n1436), .B(n1435), .Y(n865) );
  nand2a0 U1232 ( .A(n1425), .B(n1424), .Y(n870) );
  nand2a0 U1233 ( .A(n1427), .B(n1426), .Y(n869) );
  nand2a0 U1234 ( .A(n1433), .B(n1432), .Y(n866) );
  nand2a0 U1235 ( .A(n1429), .B(n1428), .Y(n868) );
  nand2a0 U1236 ( .A(n1431), .B(n1430), .Y(n867) );
  and2c0 U1237 ( .A(Instruction_27), .B(n1359), .Y(n896) );
  nand2a0 U1238 ( .A(n1356), .B(n1352), .Y(n1359) );
  and2a2 U1239 ( .A(cntrl_state_8_), .B(n972), .Y(cntrl_N106) );
  and2c0 U1240 ( .A(Reset), .B(cntrl_state_3_), .Y(n1349) );
  and2c0 U1241 ( .A(cntrl_state_1_), .B(cntrl_state_0_), .Y(n1353) );
  nand2a0 U1242 ( .A(n1387), .B(n1386), .Y(n889) );
  buf1a4 U1243 ( .A(n1439), .Y(n960) );
  nor2b2 U1244 ( .A(PCSource[0]), .B(n1437), .Y(n1438) );
  buf1a4 U1245 ( .A(n1437), .Y(n958) );
  nor2b2 U1246 ( .A(PCSource[1]), .B(n1437), .Y(n1434) );
  and2c0 U1247 ( .A(WriteAdd[0]), .B(WriteAdd[31]), .Y(n1368) );
  and2c0 U1248 ( .A(WriteAdd[2]), .B(WriteAdd[1]), .Y(n1369) );
  and2c0 U1249 ( .A(WriteAdd[4]), .B(WriteAdd[3]), .Y(n1370) );
  and2c0 U1250 ( .A(WriteAdd[8]), .B(WriteAdd[7]), .Y(n1365) );
  and2c0 U1251 ( .A(WriteAdd[10]), .B(WriteAdd[9]), .Y(n1366) );
  and2c0 U1252 ( .A(WriteAdd[22]), .B(WriteAdd[21]), .Y(n1375) );
  and2c0 U1253 ( .A(WriteAdd[24]), .B(WriteAdd[23]), .Y(n1360) );
  and2c0 U1254 ( .A(WriteAdd[28]), .B(WriteAdd[27]), .Y(n1362) );
  and2c0 U1255 ( .A(WriteAdd[30]), .B(WriteAdd[29]), .Y(n1363) );
  inv1a0 U1256 ( .A(n1442), .Y(n1444) );
  oa4f1 U1257 ( .A(MemData[8]), .B(n923), .C(n961), .D(WriteAdd[8]), .Y(n1453)
         );
  oa4f1 U1258 ( .A(MemData[0]), .B(n923), .C(n1475), .D(WriteAdd[0]), .Y(n1445) );
  inv1a0 U1259 ( .A(cntrl_state_2_), .Y(n1354) );
  and2c0 U1260 ( .A(cntrl_state_5_), .B(cntrl_state_4_), .Y(n1350) );
  inv1a0 U1261 ( .A(n1357), .Y(n1352) );
  nand2a0 U1262 ( .A(n971), .B(cntrl_state_1_), .Y(n1357) );
  and2c0 U1263 ( .A(Instruction_26), .B(Instruction_31), .Y(n1351) );
  and2c0 U1264 ( .A(Instruction_28), .B(Instruction_30), .Y(n1347) );
  oa4f1 U1265 ( .A(MemData[3]), .B(n923), .C(n1475), .D(WriteAdd[3]), .Y(n1448) );
  oa4f1 U1266 ( .A(MemData[9]), .B(n923), .C(n1475), .D(WriteAdd[9]), .Y(n1454) );
  oa4f1 U1267 ( .A(MemData[11]), .B(n962), .C(n961), .D(WriteAdd[11]), .Y(
        n1456) );
  oa4f1 U1268 ( .A(MemData[16]), .B(n923), .C(n961), .D(WriteAdd[16]), .Y(
        n1461) );
  oa4f1 U1269 ( .A(MemData[13]), .B(n962), .C(n961), .D(WriteAdd[13]), .Y(
        n1458) );
  oa4f1 U1270 ( .A(MemData[14]), .B(n962), .C(n961), .D(WriteAdd[14]), .Y(
        n1459) );
  oa4f1 U1271 ( .A(MemData[15]), .B(n923), .C(n961), .D(WriteAdd[15]), .Y(
        n1460) );
  oa4f1 U1272 ( .A(MemData[12]), .B(n923), .C(n961), .D(WriteAdd[12]), .Y(
        n1457) );
  oa4f1 U1273 ( .A(MemData[22]), .B(n962), .C(n961), .D(WriteAdd[22]), .Y(
        n1467) );
  oa4f1 U1274 ( .A(MemData[24]), .B(n923), .C(n961), .D(WriteAdd[24]), .Y(
        n1469) );
  oa4f1 U1275 ( .A(MemData[25]), .B(n962), .C(n961), .D(WriteAdd[25]), .Y(
        n1470) );
  oa4f1 U1276 ( .A(MemData[28]), .B(n962), .C(n961), .D(WriteAdd[28]), .Y(
        n1473) );
  buf1a4 U1277 ( .A(n1475), .Y(n961) );
  nor2a2 U1278 ( .A(Reset), .B(MemToReg), .Y(n1475) );
  buf1a4 U1279 ( .A(n923), .Y(n962) );
  buf1a4 U1280 ( .A(n157), .Y(n972) );
  mx2a2 U1281 ( .D0(PC[30]), .D1(WriteAdd[30]), .S(n974), .Y(ReadAdd[30]) );
  mx2a2 U1282 ( .D0(PC[29]), .D1(WriteAdd[29]), .S(IorD), .Y(ReadAdd[29]) );
  mx2a2 U1283 ( .D0(PC[28]), .D1(WriteAdd[28]), .S(IorD), .Y(ReadAdd[28]) );
  mx2a2 U1284 ( .D0(PC[27]), .D1(WriteAdd[27]), .S(n974), .Y(ReadAdd[27]) );
  mx2a2 U1285 ( .D0(PC[26]), .D1(WriteAdd[26]), .S(IorD), .Y(ReadAdd[26]) );
  mx2a2 U1286 ( .D0(PC[25]), .D1(WriteAdd[25]), .S(n974), .Y(ReadAdd[25]) );
  mx2a2 U1287 ( .D0(PC[24]), .D1(WriteAdd[24]), .S(n974), .Y(ReadAdd[24]) );
  mx2a2 U1288 ( .D0(PC[23]), .D1(WriteAdd[23]), .S(IorD), .Y(ReadAdd[23]) );
  mx2a2 U1289 ( .D0(PC[22]), .D1(WriteAdd[22]), .S(IorD), .Y(ReadAdd[22]) );
  mx2a2 U1290 ( .D0(PC[21]), .D1(WriteAdd[21]), .S(IorD), .Y(ReadAdd[21]) );
  mx2a2 U1291 ( .D0(PC[20]), .D1(WriteAdd[20]), .S(n974), .Y(ReadAdd[20]) );
  mx2a2 U1292 ( .D0(PC[19]), .D1(WriteAdd[19]), .S(IorD), .Y(ReadAdd[19]) );
  mx2a2 U1293 ( .D0(PC[18]), .D1(WriteAdd[18]), .S(n974), .Y(ReadAdd[18]) );
  mx2a2 U1294 ( .D0(PC[17]), .D1(WriteAdd[17]), .S(IorD), .Y(ReadAdd[17]) );
  mx2a2 U1295 ( .D0(PC[16]), .D1(WriteAdd[16]), .S(IorD), .Y(ReadAdd[16]) );
  mx2a2 U1296 ( .D0(PC[15]), .D1(WriteAdd[15]), .S(IorD), .Y(ReadAdd[15]) );
  mx2a2 U1297 ( .D0(PC[14]), .D1(WriteAdd[14]), .S(n974), .Y(ReadAdd[14]) );
  mx2a2 U1298 ( .D0(PC[13]), .D1(WriteAdd[13]), .S(n974), .Y(ReadAdd[13]) );
  mx2a2 U1299 ( .D0(PC[12]), .D1(WriteAdd[12]), .S(n974), .Y(ReadAdd[12]) );
  mx2a2 U1300 ( .D0(PC[11]), .D1(WriteAdd[11]), .S(n974), .Y(ReadAdd[11]) );
  mx2a2 U1301 ( .D0(PC[10]), .D1(WriteAdd[10]), .S(IorD), .Y(ReadAdd[10]) );
  mx2a2 U1302 ( .D0(PC[9]), .D1(WriteAdd[9]), .S(n974), .Y(ReadAdd[9]) );
  mx2a2 U1303 ( .D0(PC[8]), .D1(WriteAdd[8]), .S(n974), .Y(ReadAdd[8]) );
  mx2a2 U1304 ( .D0(PC[7]), .D1(WriteAdd[7]), .S(n974), .Y(ReadAdd[7]) );
  mx2a2 U1305 ( .D0(PC[6]), .D1(WriteAdd[6]), .S(n974), .Y(ReadAdd[6]) );
  mx2a2 U1306 ( .D0(PC[5]), .D1(WriteAdd[5]), .S(n974), .Y(ReadAdd[5]) );
  mx2a2 U1307 ( .D0(PC[4]), .D1(WriteAdd[4]), .S(n974), .Y(ReadAdd[4]) );
  mx2a2 U1308 ( .D0(PC[3]), .D1(WriteAdd[3]), .S(n974), .Y(ReadAdd[3]) );
  mx2a2 U1309 ( .D0(PC[2]), .D1(WriteAdd[2]), .S(n974), .Y(ReadAdd[2]) );
  mx2a2 U1310 ( .D0(PC[1]), .D1(WriteAdd[1]), .S(IorD), .Y(ReadAdd[1]) );
  mx2a2 U1311 ( .D0(PC[0]), .D1(WriteAdd[0]), .S(n974), .Y(ReadAdd[0]) );
  nand2a0 U1312 ( .A(n946), .B(alu_MuxB_30_), .Y(n1294) );
  inv1a0 U1313 ( .A(alu_MuxB_31_), .Y(n1111) );
  nand2a0 U1314 ( .A(n947), .B(alu_MuxB_29_), .Y(n1284) );
  nand2a0 U1315 ( .A(n946), .B(alu_MuxB_28_), .Y(n1280) );
  inv1a0 U1316 ( .A(alu_MuxB_29_), .Y(n1100) );
  nand2a0 U1317 ( .A(n947), .B(alu_MuxB_27_), .Y(n1276) );
  inv1a0 U1318 ( .A(alu_MuxB_28_), .Y(n1096) );
  nand2a0 U1319 ( .A(n946), .B(alu_MuxB_26_), .Y(n1272) );
  inv1a0 U1320 ( .A(alu_MuxB_27_), .Y(n1092) );
  nand2a0 U1321 ( .A(n947), .B(alu_MuxB_25_), .Y(n1268) );
  inv1a0 U1322 ( .A(alu_MuxB_26_), .Y(n1088) );
  nand2a0 U1323 ( .A(n1342), .B(alu_MuxB_24_), .Y(n1262) );
  inv1a0 U1324 ( .A(alu_MuxB_25_), .Y(n1084) );
  nand2a0 U1325 ( .A(n946), .B(alu_MuxB_23_), .Y(n1256) );
  inv1a0 U1326 ( .A(alu_MuxB_24_), .Y(n1080) );
  nand2a0 U1327 ( .A(n947), .B(alu_MuxB_22_), .Y(n1250) );
  inv1a0 U1328 ( .A(alu_MuxB_23_), .Y(n1076) );
  nand2a0 U1329 ( .A(n947), .B(alu_MuxB_21_), .Y(n1244) );
  inv1a0 U1330 ( .A(alu_MuxB_22_), .Y(n1072) );
  nand2a0 U1331 ( .A(n946), .B(alu_MuxB_20_), .Y(n1238) );
  inv1a0 U1332 ( .A(alu_MuxB_21_), .Y(n1068) );
  nand2a0 U1333 ( .A(n946), .B(alu_MuxB_19_), .Y(n1226) );
  inv1a0 U1334 ( .A(alu_MuxB_20_), .Y(n1061) );
  nand2a0 U1335 ( .A(n1342), .B(alu_MuxB_18_), .Y(n1220) );
  inv1a0 U1336 ( .A(alu_MuxB_19_), .Y(n1057) );
  nand2a0 U1337 ( .A(n947), .B(alu_MuxB_17_), .Y(n1214) );
  inv1a0 U1338 ( .A(alu_MuxB_18_), .Y(n1053) );
  nand2a0 U1339 ( .A(n946), .B(alu_MuxB_16_), .Y(n1208) );
  inv1a0 U1340 ( .A(alu_MuxB_17_), .Y(n1049) );
  mx2a2 U1341 ( .D0(PC[31]), .D1(WriteAdd[31]), .S(n974), .Y(ReadAdd[31]) );
  buf1a4 U1342 ( .A(IorD), .Y(n974) );
  nand2a0 U1343 ( .A(alu_MuxB_31_), .B(n1113), .Y(n1114) );
  nand2a0 U1344 ( .A(n948), .B(n1299), .Y(n1112) );
  and2c0 U1345 ( .A(n71), .B(n940), .Y(n1205) );
  and2c0 U1346 ( .A(n75), .B(n940), .Y(n1211) );
  and2c0 U1347 ( .A(n79), .B(n940), .Y(n1217) );
  and2c0 U1348 ( .A(n83), .B(n940), .Y(n1223) );
  and2c0 U1349 ( .A(n87), .B(n1337), .Y(n1235) );
  and2c0 U1350 ( .A(n91), .B(n940), .Y(n1241) );
  and2c0 U1351 ( .A(n95), .B(n940), .Y(n1247) );
  and2c0 U1352 ( .A(n99), .B(n940), .Y(n1253) );
  and2c0 U1353 ( .A(n103), .B(n1337), .Y(n1259) );
  and2c0 U1354 ( .A(n107), .B(n941), .Y(n1265) );
  and2c0 U1355 ( .A(n111), .B(n941), .Y(n1271) );
  and2c0 U1356 ( .A(n123), .B(n1337), .Y(n1275) );
  and2c0 U1357 ( .A(n119), .B(n940), .Y(n1279) );
  and2c0 U1358 ( .A(n115), .B(n1337), .Y(n1283) );
  and2c0 U1359 ( .A(n3), .B(n1337), .Y(n1293) );
  and2c0 U1360 ( .A(n128), .B(n1337), .Y(n1297) );
  inv1a0 U1361 ( .A(alu_MuxB_30_), .Y(n1116) );
  and2c0 U1362 ( .A(n67), .B(n940), .Y(n1199) );
  nand2a0 U1363 ( .A(n1342), .B(alu_MuxB_15_), .Y(n1202) );
  inv1a0 U1364 ( .A(alu_MuxB_16_), .Y(n1045) );
  and2c0 U1365 ( .A(n63), .B(n941), .Y(n1193) );
  nand2a0 U1366 ( .A(n947), .B(alu_MuxB_14_), .Y(n1196) );
  inv1a0 U1367 ( .A(alu_MuxB_15_), .Y(n1041) );
  and2c0 U1368 ( .A(n59), .B(n941), .Y(n1187) );
  nand2a0 U1369 ( .A(n946), .B(alu_MuxB_13_), .Y(n1190) );
  inv1a0 U1370 ( .A(alu_MuxB_12_), .Y(n1037) );
  and2c0 U1371 ( .A(n55), .B(n941), .Y(n1181) );
  nand2a0 U1372 ( .A(n946), .B(alu_MuxB_12_), .Y(n1184) );
  inv1a0 U1373 ( .A(alu_MuxB_11_), .Y(n1033) );
  and2c0 U1374 ( .A(n51), .B(n941), .Y(n1175) );
  nand2a0 U1375 ( .A(n946), .B(alu_MuxB_11_), .Y(n1178) );
  nand2a0 U1376 ( .A(n1173), .B(alu_MuxB_10_), .Y(n1024) );
  nand2a0 U1377 ( .A(n947), .B(alu_MuxA_10_), .Y(n1171) );
  and2c0 U1378 ( .A(n47), .B(n941), .Y(n1163) );
  and2c0 U1379 ( .A(n43), .B(n1337), .Y(n1341) );
  nand2a0 U1380 ( .A(n946), .B(alu_MuxB_9_), .Y(n1343) );
  inv1a0 U1381 ( .A(alu_MuxB_10_), .Y(n1147) );
  and2c0 U1382 ( .A(n39), .B(n941), .Y(n1334) );
  nand2a0 U1383 ( .A(n946), .B(alu_MuxB_8_), .Y(n1335) );
  inv1a0 U1384 ( .A(alu_MuxB_9_), .Y(n1140) );
  and2c0 U1385 ( .A(n35), .B(n941), .Y(n1324) );
  nand2a0 U1386 ( .A(n947), .B(alu_MuxB_7_), .Y(n1331) );
  inv1a0 U1387 ( .A(alu_MuxB_6_), .Y(n1136) );
  nand2a0 U1388 ( .A(n1321), .B(alu_MuxA_6_), .Y(n1127) );
  nand2a0 U1389 ( .A(n946), .B(alu_MuxB_6_), .Y(n1320) );
  nand2a0 U1390 ( .A(n1322), .B(alu_MuxB_6_), .Y(n1128) );
  nand2a0 U1391 ( .A(n1132), .B(alu_MuxB_7_), .Y(n1129) );
  and2c0 U1392 ( .A(n31), .B(n940), .Y(n1317) );
  and2c0 U1393 ( .A(n27), .B(n1337), .Y(n1313) );
  nand2a0 U1394 ( .A(n1311), .B(alu_MuxA_4_), .Y(n1122) );
  nand2a0 U1395 ( .A(n946), .B(alu_MuxB_4_), .Y(n1310) );
  nand2a0 U1396 ( .A(n1143), .B(alu_MuxB_3_), .Y(n1123) );
  inv1a4 U1397 ( .A(n1135), .Y(n1143) );
  nand2a0 U1398 ( .A(alu_MuxB_4_), .B(n1121), .Y(n1124) );
  and2c0 U1399 ( .A(n23), .B(n941), .Y(n1307) );
  and2c0 U1400 ( .A(n19), .B(n1337), .Y(n1301) );
  nand2a0 U1401 ( .A(n947), .B(alu_MuxB_3_), .Y(n1304) );
  inv1a0 U1402 ( .A(alu_MuxB_2_), .Y(n1120) );
  and2c0 U1403 ( .A(n15), .B(n941), .Y(n1287) );
  inv1a0 U1404 ( .A(WriteData[2]), .Y(n1014) );
  and2c0 U1405 ( .A(n11), .B(n940), .Y(n1229) );
  or2c2 U1406 ( .A(n1023), .B(n1022), .Y(n1135) );
  nand2a0 U1407 ( .A(n924), .B(n1019), .Y(n1020) );
  or3b2 U1408 ( .B(n1018), .C(ALUOp[0]), .A(ALUOp[1]), .Y(n1141) );
  inv1a0 U1409 ( .A(n1159), .Y(n1017) );
  nand2a0 U1410 ( .A(Read1RegSel[0]), .B(n1154), .Y(n1338) );
  and2c0 U1411 ( .A(n7), .B(n941), .Y(n1156) );
  buf1a4 U1412 ( .A(n1011), .Y(n928) );
  and2c0 U1413 ( .A(n973), .B(Read1RegSel[1]), .Y(n1154) );
  buf1a4 U1414 ( .A(n139), .Y(n973) );
  nand2a0 U1415 ( .A(n924), .B(n947), .Y(n1160) );
  and2c0 U1416 ( .A(n1149), .B(n1170), .Y(n1342) );
  inv1a2 U1417 ( .A(n930), .Y(n929) );
  inv1a4 U1418 ( .A(n1132), .Y(n1146) );
  nor2a2 U1419 ( .A(Instruction[5]), .B(n1159), .Y(n1132) );
  inv1a0 U1420 ( .A(alu_MuxB_1_), .Y(n1107) );
  nor2a2 U1421 ( .A(ALUSelB[1]), .B(ALUSelB[0]), .Y(n1013) );
  inv1a0 U1422 ( .A(WriteData[1]), .Y(n1016) );
  nand2a0 U1423 ( .A(n1150), .B(n1151), .Y(n1326) );
  or2c2 U1424 ( .A(Read2RegSel[1]), .B(n1150), .Y(n1330) );
  mx2d0 U1425 ( .D0(n1455), .D1(n48), .S(n970), .Y(n819) );
  buf1a2 U1426 ( .A(n970), .Y(n969) );
  mx2d0 U1427 ( .D0(n1455), .D1(n46), .S(n968), .Y(n821) );
  buf1a2 U1428 ( .A(n968), .Y(n967) );
  buf1a2 U1429 ( .A(n965), .Y(n966) );
  oa1d1 U1430 ( .A(n1440), .B(n1444), .C(Reset), .Y(n1478) );
  or4e0 U1431 ( .A(n1347), .B(Instruction_26), .C(Instruction_31), .D(
        Instruction_27), .Y(n1358) );
  buf1a2 U1432 ( .A(n963), .Y(n964) );
  oa1d1 U1433 ( .A(n1442), .B(n1440), .C(Reset), .Y(n1476) );
  buf1a2 U1434 ( .A(n972), .Y(n971) );
  buf1a2 U1435 ( .A(n1344), .Y(n951) );
  nand2a0 U1436 ( .A(Read2RegSel[0]), .B(n1151), .Y(n1325) );
  buf1a2 U1437 ( .A(n1328), .Y(n937) );
  buf1a2 U1438 ( .A(n939), .Y(n938) );
  ao1d1 U1439 ( .A(n929), .B(WriteData[17]), .C(n1012), .Y(alu_MuxB_17_) );
  ao1d1 U1440 ( .A(n1013), .B(WriteData[18]), .C(n1012), .Y(alu_MuxB_18_) );
  ao1d1 U1441 ( .A(n1013), .B(WriteData[19]), .C(n1012), .Y(alu_MuxB_19_) );
  ao1d1 U1442 ( .A(n1013), .B(WriteData[20]), .C(n1012), .Y(alu_MuxB_20_) );
  ao1d1 U1443 ( .A(n929), .B(WriteData[21]), .C(n1012), .Y(alu_MuxB_21_) );
  ao1d1 U1444 ( .A(n1013), .B(WriteData[22]), .C(n1012), .Y(alu_MuxB_22_) );
  ao1d1 U1445 ( .A(n1013), .B(WriteData[23]), .C(n1012), .Y(alu_MuxB_23_) );
  ao1d1 U1446 ( .A(n1013), .B(WriteData[24]), .C(n1012), .Y(alu_MuxB_24_) );
  ao1d1 U1447 ( .A(n1013), .B(WriteData[25]), .C(n925), .Y(alu_MuxB_25_) );
  ao1d1 U1448 ( .A(n929), .B(WriteData[26]), .C(n925), .Y(alu_MuxB_26_) );
  ao1d1 U1449 ( .A(n929), .B(WriteData[27]), .C(n925), .Y(alu_MuxB_27_) );
  ao1d1 U1450 ( .A(n929), .B(WriteData[28]), .C(n925), .Y(alu_MuxB_28_) );
  ao1d1 U1451 ( .A(n929), .B(WriteData[29]), .C(n925), .Y(alu_MuxB_29_) );
  ao1d1 U1452 ( .A(n929), .B(WriteData[31]), .C(n925), .Y(alu_MuxB_31_) );
  ao1d1 U1453 ( .A(n929), .B(WriteData[30]), .C(n925), .Y(alu_MuxB_30_) );
  ao1d1 U1454 ( .A(n1013), .B(WriteData[16]), .C(n925), .Y(alu_MuxB_16_) );
  ao1d1 U1455 ( .A(n1013), .B(WriteData[15]), .C(n925), .Y(alu_MuxB_15_) );
  ao1f1 U1456 ( .A(n938), .B(n7), .C(n1153), .Y(WriteData[0]) );
  ao1f1 U1457 ( .A(n938), .B(n111), .C(n1267), .Y(WriteData[26]) );
  ao1f1 U1458 ( .A(n1330), .B(n107), .C(n1261), .Y(WriteData[25]) );
  ao1f1 U1459 ( .A(n939), .B(n103), .C(n1255), .Y(WriteData[24]) );
  ao1f1 U1460 ( .A(n938), .B(n95), .C(n1243), .Y(WriteData[22]) );
  ao1f1 U1461 ( .A(n939), .B(n83), .C(n1219), .Y(WriteData[19]) );
  ao1f1 U1462 ( .A(n939), .B(n79), .C(n1213), .Y(WriteData[18]) );
  ao1f1 U1463 ( .A(n939), .B(n75), .C(n1207), .Y(WriteData[17]) );
  ao1f1 U1464 ( .A(n939), .B(n55), .C(n1177), .Y(WriteData[12]) );
  ao1f1 U1465 ( .A(n47), .B(n1330), .C(n1169), .Y(WriteData[10]) );
  ao1f1 U1466 ( .A(n939), .B(n43), .C(n1165), .Y(WriteData[9]) );
  ao1f1 U1467 ( .A(n938), .B(n35), .C(n1319), .Y(WriteData[7]) );
  ao1f1 U1468 ( .A(n938), .B(n31), .C(n1315), .Y(WriteData[6]) );
  ao1f1 U1469 ( .A(n27), .B(n939), .C(n1309), .Y(WriteData[5]) );
  ao1f1 U1470 ( .A(n938), .B(n15), .C(n1231), .Y(WriteData[2]) );
  ao1f1 U1471 ( .A(n938), .B(n11), .C(n1158), .Y(WriteData[1]) );
  or4a1 U1472 ( .A(n1355), .B(cntrl_N114), .C(cntrl_N111), .D(n155), .Y(
        cntrl_N113) );
  nor2b1 U1473 ( .A(n155), .B(n419), .Y(cntrl_N103) );
  nor2a1 U1474 ( .A(Instruction_29), .B(n1358), .Y(n419) );
  ao7a2 U1475 ( .A(WriteAdd[31]), .B(n960), .C(n1438), .D(TargetReg[31]), .E(
        PC[31]), .F(n958), .Y(n863) );
  ao7a2 U1476 ( .A(WriteAdd[30]), .B(n1439), .C(n959), .D(TargetReg[30]), .E(
        PC[30]), .F(n1437), .Y(n864) );
  or4e0 U1477 ( .A(n1350), .B(n1353), .C(n1349), .D(n1354), .Y(cntrl_N109) );
  or4e0 U1478 ( .A(n1375), .B(n1374), .C(n1373), .D(n1372), .Y(n1376) );
  or4e0 U1479 ( .A(n1370), .B(n1369), .C(PCWriteCond), .D(n1368), .Y(n1371) );
  or4c0 U1480 ( .C(WriteAdd[12]), .D(WriteAdd[11]), .A(n1366), .B(n1365), .Y(
        n1367) );
  or4a1 U1481 ( .A(WriteAdd[18]), .B(WriteAdd[17]), .C(WriteAdd[16]), .D(
        WriteAdd[15]), .Y(n1364) );
  or4e0 U1482 ( .A(n1363), .B(n1362), .C(n1361), .D(n1360), .Y(n1377) );
  or3b1 U1483 ( .B(cntrl_state_9_), .C(cntrl_state_10_), .A(n1350), .Y(n426)
         );
  nor3c1 U1484 ( .A(n1352), .B(n1358), .C(n145), .Y(n1355) );
  nor3c1 U1485 ( .A(n1347), .B(n1351), .C(Instruction_29), .Y(n1356) );
  oa4f0 U1486 ( .A(n1143), .B(alu_MuxB_29_), .C(alu_MuxB_30_), .D(n1108), .Y(
        n1109) );
  oa4f0 U1487 ( .A(n1295), .B(alu_MuxA_30_), .C(C55_DATA6_30), .D(n931), .Y(
        n1110) );
  oa4f0 U1488 ( .A(n1143), .B(alu_MuxB_28_), .C(alu_MuxB_29_), .D(n1101), .Y(
        n1102) );
  oa4f0 U1489 ( .A(n1285), .B(alu_MuxA_29_), .C(C55_DATA6_29), .D(n1141), .Y(
        n1103) );
  oa4f0 U1490 ( .A(n1143), .B(alu_MuxB_27_), .C(alu_MuxB_28_), .D(n1097), .Y(
        n1098) );
  oa4f0 U1491 ( .A(n1281), .B(alu_MuxA_28_), .C(C55_DATA6_28), .D(n1141), .Y(
        n1099) );
  oa4f0 U1492 ( .A(n1143), .B(alu_MuxB_26_), .C(alu_MuxB_27_), .D(n1093), .Y(
        n1094) );
  oa4f0 U1493 ( .A(n1277), .B(alu_MuxA_27_), .C(C55_DATA6_27), .D(n931), .Y(
        n1095) );
  oa4f0 U1494 ( .A(n1143), .B(alu_MuxB_25_), .C(alu_MuxB_26_), .D(n1089), .Y(
        n1090) );
  oa4f0 U1495 ( .A(n1273), .B(alu_MuxA_26_), .C(C55_DATA6_26), .D(n1141), .Y(
        n1091) );
  oa4f0 U1496 ( .A(n1143), .B(alu_MuxB_24_), .C(alu_MuxB_25_), .D(n1085), .Y(
        n1086) );
  oa4f0 U1497 ( .A(n1269), .B(alu_MuxA_25_), .C(C55_DATA6_25), .D(n1141), .Y(
        n1087) );
  oa4f0 U1498 ( .A(n1143), .B(alu_MuxB_23_), .C(alu_MuxB_24_), .D(n1081), .Y(
        n1082) );
  oa4f0 U1499 ( .A(n1263), .B(alu_MuxA_24_), .C(C55_DATA6_24), .D(n1141), .Y(
        n1083) );
  oa4f0 U1500 ( .A(n1143), .B(alu_MuxB_22_), .C(alu_MuxB_23_), .D(n1077), .Y(
        n1078) );
  oa4f0 U1501 ( .A(n1257), .B(alu_MuxA_23_), .C(C55_DATA6_23), .D(n1141), .Y(
        n1079) );
  oa4f0 U1502 ( .A(n1143), .B(alu_MuxB_21_), .C(alu_MuxB_22_), .D(n1073), .Y(
        n1074) );
  oa4f0 U1503 ( .A(n1251), .B(alu_MuxA_22_), .C(C55_DATA6_22), .D(n931), .Y(
        n1075) );
  oa4f0 U1504 ( .A(n1143), .B(alu_MuxB_20_), .C(alu_MuxB_21_), .D(n1069), .Y(
        n1070) );
  oa4f0 U1505 ( .A(n1245), .B(alu_MuxA_21_), .C(C55_DATA6_21), .D(n1141), .Y(
        n1071) );
  oa4f0 U1506 ( .A(n1143), .B(alu_MuxB_19_), .C(alu_MuxB_20_), .D(n1065), .Y(
        n1066) );
  oa4f0 U1507 ( .A(n1239), .B(alu_MuxA_20_), .C(C55_DATA6_20), .D(n931), .Y(
        n1067) );
  oa4f0 U1508 ( .A(n1143), .B(alu_MuxB_18_), .C(alu_MuxB_19_), .D(n1058), .Y(
        n1059) );
  oa4f0 U1509 ( .A(n1227), .B(alu_MuxA_19_), .C(C55_DATA6_19), .D(n931), .Y(
        n1060) );
  oa4f0 U1510 ( .A(n1143), .B(alu_MuxB_17_), .C(alu_MuxB_18_), .D(n1054), .Y(
        n1055) );
  oa4f0 U1511 ( .A(n1221), .B(alu_MuxA_18_), .C(C55_DATA6_18), .D(n931), .Y(
        n1056) );
  oa4f0 U1512 ( .A(n1143), .B(alu_MuxB_16_), .C(alu_MuxB_17_), .D(n1050), .Y(
        n1051) );
  oa4f0 U1513 ( .A(n1215), .B(alu_MuxA_17_), .C(C55_DATA6_17), .D(n931), .Y(
        n1052) );
  oa4f0 U1514 ( .A(n1143), .B(alu_MuxB_15_), .C(alu_MuxB_16_), .D(n1046), .Y(
        n1047) );
  oa4f0 U1515 ( .A(n1209), .B(alu_MuxA_16_), .C(C55_DATA6_16), .D(n931), .Y(
        n1048) );
  oa4f0 U1516 ( .A(C55_DATA6_31), .B(n1141), .C(alu_MuxA_31_), .D(n1112), .Y(
        n1115) );
  oa2i0 U1517 ( .A(PC[16]), .B(n973), .C(n1205), .D(n1204), .Y(n995) );
  oa2i0 U1518 ( .A(PC[17]), .B(n139), .C(n1211), .D(n1210), .Y(n994) );
  oa2i0 U1519 ( .A(PC[18]), .B(n139), .C(n1217), .D(n1216), .Y(n993) );
  oa2i0 U1520 ( .A(PC[19]), .B(n973), .C(n1223), .D(n1222), .Y(n992) );
  oa2i0 U1521 ( .A(PC[20]), .B(n973), .C(n1235), .D(n1234), .Y(n991) );
  oa2i0 U1522 ( .A(PC[21]), .B(n139), .C(n1241), .D(n1240), .Y(n990) );
  oa2i0 U1523 ( .A(PC[22]), .B(n139), .C(n1247), .D(n1246), .Y(n989) );
  oa2i0 U1524 ( .A(PC[23]), .B(n973), .C(n1253), .D(n1252), .Y(n988) );
  oa2i0 U1525 ( .A(PC[24]), .B(n973), .C(n1259), .D(n1258), .Y(n987) );
  oa2i0 U1526 ( .A(PC[25]), .B(n139), .C(n1265), .D(n1264), .Y(n986) );
  oa2i0 U1527 ( .A(PC[26]), .B(n973), .C(n1271), .D(n1270), .Y(n985) );
  oa2i0 U1528 ( .A(PC[27]), .B(n139), .C(n1275), .D(n1274), .Y(n984) );
  oa2i0 U1529 ( .A(PC[28]), .B(n973), .C(n1279), .D(n1278), .Y(n983) );
  oa2i0 U1530 ( .A(PC[29]), .B(n973), .C(n1283), .D(n1282), .Y(n982) );
  oa2i0 U1531 ( .A(PC[30]), .B(n973), .C(n1293), .D(n1292), .Y(n981) );
  oa2i0 U1532 ( .A(PC[31]), .B(n139), .C(n1297), .D(n1296), .Y(n980) );
  oa4f0 U1533 ( .A(n1143), .B(alu_MuxB_14_), .C(alu_MuxB_15_), .D(n1042), .Y(
        n1043) );
  oa4f0 U1534 ( .A(n1203), .B(alu_MuxA_15_), .C(C55_DATA6_15), .D(n931), .Y(
        n1044) );
  oa2i0 U1535 ( .A(PC[15]), .B(n139), .C(n1199), .D(n1198), .Y(n996) );
  oa4f0 U1536 ( .A(n1143), .B(alu_MuxB_13_), .C(alu_MuxB_14_), .D(n1038), .Y(
        n1039) );
  oa4f0 U1537 ( .A(n1197), .B(alu_MuxA_14_), .C(C55_DATA6_14), .D(n931), .Y(
        n1040) );
  oa2i0 U1538 ( .A(PC[14]), .B(n973), .C(n1193), .D(n1192), .Y(n997) );
  oa4f0 U1539 ( .A(n1132), .B(alu_MuxB_14_), .C(alu_MuxB_13_), .D(n1034), .Y(
        n1035) );
  ao4a2 U1540 ( .A(n929), .B(WriteData[14]), .C(ALUSelB[1]), .D(
        Instruction[14]), .Y(alu_MuxB_14_) );
  oa4f0 U1541 ( .A(n1191), .B(alu_MuxA_13_), .C(C55_DATA6_13), .D(n931), .Y(
        n1036) );
  oa2i0 U1542 ( .A(PC[13]), .B(n139), .C(n1187), .D(n1186), .Y(n998) );
  oa4f0 U1543 ( .A(n1132), .B(alu_MuxB_13_), .C(alu_MuxB_12_), .D(n1030), .Y(
        n1031) );
  ao4a2 U1544 ( .A(n1013), .B(WriteData[13]), .C(ALUSelB[1]), .D(
        Instruction[13]), .Y(alu_MuxB_13_) );
  oa4f0 U1545 ( .A(n1185), .B(alu_MuxA_12_), .C(C55_DATA6_12), .D(n1141), .Y(
        n1032) );
  oa2i0 U1546 ( .A(PC[12]), .B(n973), .C(n1181), .D(n1180), .Y(n999) );
  oa4f0 U1547 ( .A(n1132), .B(alu_MuxB_12_), .C(alu_MuxB_11_), .D(n1027), .Y(
        n1028) );
  ao4a2 U1548 ( .A(n929), .B(WriteData[12]), .C(ALUSelB[1]), .D(
        Instruction[12]), .Y(alu_MuxB_12_) );
  oa4f0 U1549 ( .A(n1179), .B(alu_MuxA_11_), .C(C55_DATA6_11), .D(n931), .Y(
        n1029) );
  oa2i0 U1550 ( .A(PC[11]), .B(n973), .C(n1175), .D(n1174), .Y(n1000) );
  oa4f0 U1551 ( .A(n1143), .B(alu_MuxB_9_), .C(n1132), .D(alu_MuxB_11_), .Y(
        n1025) );
  ao4a2 U1552 ( .A(n1013), .B(WriteData[11]), .C(ALUSelB[1]), .D(
        Instruction[11]), .Y(alu_MuxB_11_) );
  oa4f0 U1553 ( .A(n1172), .B(alu_MuxA_10_), .C(C55_DATA6_10), .D(n931), .Y(
        n1026) );
  oa2i0 U1554 ( .A(PC[10]), .B(n139), .C(n1163), .D(n1162), .Y(n1001) );
  oa4f0 U1555 ( .A(n1143), .B(alu_MuxB_8_), .C(alu_MuxB_9_), .D(n1142), .Y(
        n1144) );
  oa4f0 U1556 ( .A(n1346), .B(alu_MuxA_9_), .C(C55_DATA6_9), .D(n931), .Y(
        n1145) );
  oa2i0 U1557 ( .A(PC[9]), .B(n973), .C(n1341), .D(n1340), .Y(n1002) );
  ao4a2 U1558 ( .A(Instruction[10]), .B(ALUSelB[1]), .C(n929), .D(
        WriteData[10]), .Y(alu_MuxB_10_) );
  oa4f0 U1559 ( .A(n1143), .B(alu_MuxB_7_), .C(alu_MuxB_8_), .D(n1137), .Y(
        n1138) );
  oa4f0 U1560 ( .A(n1336), .B(alu_MuxA_8_), .C(C55_DATA6_8), .D(n1141), .Y(
        n1139) );
  oa2i0 U1561 ( .A(PC[8]), .B(n139), .C(n1334), .D(n1333), .Y(n1003) );
  ao4a2 U1562 ( .A(n929), .B(WriteData[9]), .C(ALUSelB[1]), .D(Instruction[9]), 
        .Y(alu_MuxB_9_) );
  oa4f0 U1563 ( .A(n1132), .B(alu_MuxB_8_), .C(alu_MuxB_7_), .D(n1131), .Y(
        n1133) );
  ao4a2 U1564 ( .A(n929), .B(WriteData[8]), .C(ALUSelB[1]), .D(Instruction[8]), 
        .Y(alu_MuxB_8_) );
  oa4f0 U1565 ( .A(n1332), .B(alu_MuxA_7_), .C(C55_DATA6_7), .D(n1141), .Y(
        n1134) );
  oa2i0 U1566 ( .A(PC[7]), .B(n139), .C(n1324), .D(n1323), .Y(n1004) );
  ao4a2 U1567 ( .A(n929), .B(WriteData[7]), .C(ALUSelB[1]), .D(Instruction[7]), 
        .Y(alu_MuxB_7_) );
  oa4f0 U1568 ( .A(n1143), .B(n1126), .C(C55_DATA6_6), .D(n1141), .Y(n1130) );
  oa2i0 U1569 ( .A(PC[6]), .B(n139), .C(n1317), .D(n1316), .Y(n1005) );
  ao4a2 U1570 ( .A(n1013), .B(WriteData[6]), .C(ALUSelB[1]), .D(Instruction[6]), .Y(alu_MuxB_6_) );
  oa2i0 U1571 ( .A(PC[5]), .B(n973), .C(n1313), .D(n1312), .Y(n1006) );
  oa4f0 U1572 ( .A(n1126), .B(n1132), .C(C55_DATA6_4), .D(n1141), .Y(n1125) );
  oa2i0 U1573 ( .A(PC[4]), .B(n973), .C(n1307), .D(n1306), .Y(n1007) );
  oa4f0 U1574 ( .A(n1132), .B(alu_MuxB_4_), .C(alu_MuxB_3_), .D(n1117), .Y(
        n1118) );
  ao4a2 U1575 ( .A(n929), .B(WriteData[4]), .C(ALUSelB[1]), .D(Instruction[4]), 
        .Y(alu_MuxB_4_) );
  oa4f0 U1576 ( .A(n1305), .B(alu_MuxA_3_), .C(C55_DATA6_3), .D(n1141), .Y(
        n1119) );
  oa2i0 U1577 ( .A(PC[3]), .B(n973), .C(n1301), .D(n1300), .Y(n1008) );
  oa4f0 U1578 ( .A(n1132), .B(alu_MuxB_3_), .C(alu_MuxB_2_), .D(n1104), .Y(
        n1105) );
  ao4a2 U1579 ( .A(n1013), .B(WriteData[3]), .C(ALUSelB[1]), .D(Instruction[3]), .Y(alu_MuxB_3_) );
  oa4f0 U1580 ( .A(n1291), .B(alu_MuxA_2_), .C(C55_DATA6_2), .D(n931), .Y(
        n1106) );
  oa2i0 U1581 ( .A(PC[2]), .B(n139), .C(n1287), .D(n1286), .Y(n1009) );
  oa4f0 U1582 ( .A(n1132), .B(alu_MuxB_2_), .C(alu_MuxB_1_), .D(n1062), .Y(
        n1063) );
  oa4f0 U1583 ( .A(n1233), .B(alu_MuxA_1_), .C(C55_DATA6_1), .D(n1141), .Y(
        n1064) );
  oa2i0 U1584 ( .A(PC[1]), .B(n139), .C(n1229), .D(n1228), .Y(n1010) );
  inv1a1 U1585 ( .A(n1170), .Y(n1023) );
  oa4f0 U1586 ( .A(n1161), .B(alu_MuxA_0_), .C(C55_DATA6_0), .D(n931), .Y(
        n1021) );
  oa2i0 U1587 ( .A(PC[0]), .B(n139), .C(n1156), .D(n1155), .Y(n979) );
  or3b1 U1588 ( .B(Read1RegSel[0]), .C(n973), .A(Read1RegSel[1]), .Y(n1337) );
  inv1a1 U1589 ( .A(ALUSelB[1]), .Y(n1015) );
  buf1a2 U1590 ( .A(n1339), .Y(n945) );
  buf1a2 U1591 ( .A(n1326), .Y(n935) );
  buf1a2 U1592 ( .A(n1338), .Y(n942) );
  buf1a2 U1593 ( .A(n1325), .Y(n933) );
  buf1a2 U1594 ( .A(n1342), .Y(n947) );
  buf1a2 U1595 ( .A(n951), .Y(n948) );
  buf1a2 U1596 ( .A(n951), .Y(n950) );
  buf1a2 U1597 ( .A(n1326), .Y(n934) );
  buf1a2 U1598 ( .A(n1339), .Y(n944) );
  buf1a2 U1599 ( .A(n942), .Y(n943) );
  buf1a2 U1600 ( .A(n1325), .Y(n932) );
  buf1a2 U1601 ( .A(IRWrite), .Y(n978) );
  buf1a2 U1602 ( .A(IRWrite), .Y(n977) );
  buf1a2 U1603 ( .A(TargetWrite), .Y(n976) );
  buf1a2 U1604 ( .A(TargetWrite), .Y(n975) );
  buf1a2 U1605 ( .A(n1141), .Y(n931) );
  buf1a2 U1606 ( .A(n1345), .Y(n955) );
  buf1a2 U1607 ( .A(n1345), .Y(n954) );
  buf1a2 U1608 ( .A(n1345), .Y(n953) );
  buf1a2 U1609 ( .A(n1345), .Y(n952) );
  buf1a2 U1610 ( .A(n1337), .Y(n940) );
  buf1a2 U1611 ( .A(n1337), .Y(n941) );
  buf1a2 U1612 ( .A(n937), .Y(n936) );
  buf1a2 U1613 ( .A(n947), .Y(n946) );
  vdd U1614 ( .Y(n144) );
  gnd U1615 ( .Y(n142) );
  buf1a2 U1616 ( .A(DP_OP_100J1_124_3689_n100), .Y(n926) );
  buf1a2 U1617 ( .A(DP_OP_100J1_124_3689_n100), .Y(n927) );
  ao1f1 U1618 ( .A(n5), .B(n928), .C(n979), .Y(alu_MuxA_0_) );
  ao1f1 U1619 ( .A(n125), .B(n928), .C(n980), .Y(alu_MuxA_31_) );
  ao1f1 U1620 ( .A(n1), .B(n928), .C(n981), .Y(alu_MuxA_30_) );
  ao1f1 U1621 ( .A(n113), .B(n928), .C(n982), .Y(alu_MuxA_29_) );
  ao1f1 U1622 ( .A(n117), .B(n928), .C(n983), .Y(alu_MuxA_28_) );
  ao1f1 U1623 ( .A(n121), .B(n928), .C(n984), .Y(alu_MuxA_27_) );
  ao1f1 U1624 ( .A(n109), .B(n928), .C(n985), .Y(alu_MuxA_26_) );
  ao1f1 U1625 ( .A(n105), .B(n928), .C(n986), .Y(alu_MuxA_25_) );
  ao1f1 U1626 ( .A(n101), .B(n1011), .C(n987), .Y(alu_MuxA_24_) );
  ao1f1 U1627 ( .A(n97), .B(n928), .C(n988), .Y(alu_MuxA_23_) );
  ao1f1 U1628 ( .A(n93), .B(n928), .C(n989), .Y(alu_MuxA_22_) );
  ao1f1 U1629 ( .A(n89), .B(n928), .C(n990), .Y(alu_MuxA_21_) );
  ao1f1 U1630 ( .A(n85), .B(n928), .C(n991), .Y(alu_MuxA_20_) );
  ao1f1 U1631 ( .A(n81), .B(n928), .C(n992), .Y(alu_MuxA_19_) );
  ao1f1 U1632 ( .A(n77), .B(n928), .C(n993), .Y(alu_MuxA_18_) );
  ao1f1 U1633 ( .A(n73), .B(n928), .C(n994), .Y(alu_MuxA_17_) );
  ao1f1 U1634 ( .A(n69), .B(n928), .C(n995), .Y(alu_MuxA_16_) );
  ao1f1 U1635 ( .A(n65), .B(n928), .C(n996), .Y(alu_MuxA_15_) );
  ao1f1 U1636 ( .A(n61), .B(n1011), .C(n997), .Y(alu_MuxA_14_) );
  ao1f1 U1637 ( .A(n57), .B(n928), .C(n998), .Y(alu_MuxA_13_) );
  ao1f1 U1638 ( .A(n53), .B(n1011), .C(n999), .Y(alu_MuxA_12_) );
  ao1f1 U1639 ( .A(n49), .B(n1011), .C(n1000), .Y(alu_MuxA_11_) );
  ao1f1 U1640 ( .A(n45), .B(n928), .C(n1001), .Y(alu_MuxA_10_) );
  ao1f1 U1641 ( .A(n41), .B(n928), .C(n1002), .Y(alu_MuxA_9_) );
  ao1f1 U1642 ( .A(n37), .B(n1011), .C(n1003), .Y(alu_MuxA_8_) );
  ao1f1 U1643 ( .A(n33), .B(n928), .C(n1004), .Y(alu_MuxA_7_) );
  ao1f1 U1644 ( .A(n29), .B(n928), .C(n1005), .Y(alu_MuxA_6_) );
  ao1f1 U1645 ( .A(n25), .B(n1011), .C(n1006), .Y(alu_MuxA_5_) );
  ao1f1 U1646 ( .A(n21), .B(n928), .C(n1007), .Y(alu_MuxA_4_) );
  ao1f1 U1647 ( .A(n17), .B(n928), .C(n1008), .Y(alu_MuxA_3_) );
  ao1f1 U1648 ( .A(n13), .B(n1011), .C(n1009), .Y(alu_MuxA_2_) );
  ao1f1 U1649 ( .A(n9), .B(n1011), .C(n1010), .Y(alu_MuxA_1_) );
  ao1f1 U1650 ( .A(n938), .B(n71), .C(n1201), .Y(WriteData[16]) );
  ao1f1 U1651 ( .A(n1330), .B(n67), .C(n1195), .Y(WriteData[15]) );
  ao1f1 U1652 ( .A(n939), .B(n63), .C(n1189), .Y(WriteData[14]) );
  ao1f1 U1653 ( .A(n939), .B(n59), .C(n1183), .Y(WriteData[13]) );
  ao1f1 U1654 ( .A(n938), .B(n51), .C(n1167), .Y(WriteData[11]) );
  ao1f1 U1655 ( .A(n939), .B(n39), .C(n1329), .Y(WriteData[8]) );
  ao1f1 U1656 ( .A(n938), .B(n23), .C(n1303), .Y(WriteData[4]) );
  ao1f1 U1657 ( .A(n938), .B(n19), .C(n1289), .Y(WriteData[3]) );
  ao1f1 U1658 ( .A(n1345), .B(alu_MuxA_0_), .C(n950), .Y(n1019) );
  ao1f1 U1659 ( .A(alu_MuxA_11_), .B(n955), .C(n948), .Y(n1027) );
  ao1f1 U1660 ( .A(n953), .B(alu_MuxA_12_), .C(n951), .Y(n1030) );
  ao1f1 U1661 ( .A(n954), .B(alu_MuxA_13_), .C(n950), .Y(n1034) );
  ao1f1 U1662 ( .A(n955), .B(alu_MuxA_14_), .C(n951), .Y(n1038) );
  ao1f1 U1663 ( .A(n955), .B(alu_MuxA_15_), .C(n948), .Y(n1042) );
  ao1f1 U1664 ( .A(n953), .B(alu_MuxA_16_), .C(n948), .Y(n1046) );
  ao1f1 U1665 ( .A(n954), .B(alu_MuxA_17_), .C(n951), .Y(n1050) );
  ao1f1 U1666 ( .A(n955), .B(alu_MuxA_18_), .C(n948), .Y(n1054) );
  ao1f1 U1667 ( .A(n1345), .B(alu_MuxA_19_), .C(n951), .Y(n1058) );
  ao1f1 U1668 ( .A(n952), .B(alu_MuxA_1_), .C(n951), .Y(n1062) );
  ao1f1 U1669 ( .A(n1345), .B(alu_MuxA_20_), .C(n951), .Y(n1065) );
  ao1f1 U1670 ( .A(n1345), .B(alu_MuxA_21_), .C(n951), .Y(n1069) );
  ao1f1 U1671 ( .A(n955), .B(alu_MuxA_22_), .C(n951), .Y(n1073) );
  ao1f1 U1672 ( .A(n955), .B(alu_MuxA_23_), .C(n948), .Y(n1077) );
  ao1f1 U1673 ( .A(n954), .B(alu_MuxA_24_), .C(n951), .Y(n1081) );
  ao1f1 U1674 ( .A(n952), .B(alu_MuxA_25_), .C(n950), .Y(n1085) );
  ao1f1 U1675 ( .A(n952), .B(alu_MuxA_26_), .C(n950), .Y(n1089) );
  ao1f1 U1676 ( .A(n1345), .B(alu_MuxA_27_), .C(n949), .Y(n1093) );
  ao1f1 U1677 ( .A(n1345), .B(alu_MuxA_28_), .C(n949), .Y(n1097) );
  ao1f1 U1678 ( .A(n954), .B(alu_MuxA_29_), .C(n949), .Y(n1101) );
  ao1f1 U1679 ( .A(n954), .B(alu_MuxA_2_), .C(n949), .Y(n1104) );
  ao1f1 U1680 ( .A(n952), .B(alu_MuxA_30_), .C(n949), .Y(n1108) );
  ao1f1 U1681 ( .A(n953), .B(alu_MuxA_31_), .C(n950), .Y(n1113) );
  ao1f1 U1682 ( .A(n952), .B(alu_MuxA_3_), .C(n949), .Y(n1117) );
  ao1f1 U1683 ( .A(n953), .B(alu_MuxA_4_), .C(n948), .Y(n1121) );
  ao1f1 U1684 ( .A(n954), .B(alu_MuxA_7_), .C(n948), .Y(n1131) );
  ao1f1 U1685 ( .A(n955), .B(alu_MuxA_8_), .C(n948), .Y(n1137) );
  ao1f1 U1686 ( .A(n955), .B(alu_MuxA_9_), .C(n948), .Y(n1142) );
  ao4f0 U1687 ( .A(n5), .B(n934), .C(n6), .D(n932), .Y(n1152) );
  oa1d1 U1688 ( .A(n8), .B(n936), .C(n1152), .Y(n1153) );
  ao4f0 U1689 ( .A(n6), .B(n942), .C(n8), .D(n1339), .Y(n1155) );
  ao4f0 U1690 ( .A(n9), .B(n934), .C(n10), .D(n932), .Y(n1157) );
  oa1d1 U1691 ( .A(n12), .B(n937), .C(n1157), .Y(n1158) );
  ao2i0 U1692 ( .A(n953), .B(n924), .C(n950), .D(n1160), .Y(n1161) );
  ao4f0 U1693 ( .A(n48), .B(n945), .C(n46), .D(n943), .Y(n1162) );
  ao4f0 U1694 ( .A(n41), .B(n935), .C(n42), .D(n932), .Y(n1164) );
  oa1d1 U1695 ( .A(n44), .B(n1328), .C(n1164), .Y(n1165) );
  ao4f0 U1696 ( .A(n49), .B(n935), .C(n50), .D(n932), .Y(n1166) );
  oa1d1 U1697 ( .A(n52), .B(n937), .C(n1166), .Y(n1167) );
  ao4f0 U1698 ( .A(n45), .B(n934), .C(n46), .D(n932), .Y(n1168) );
  oa1d1 U1699 ( .A(n48), .B(n936), .C(n1168), .Y(n1169) );
  ao2i0 U1700 ( .A(n952), .B(alu_MuxA_10_), .C(n950), .D(n1171), .Y(n1173) );
  ao1f1 U1701 ( .A(n953), .B(alu_MuxB_10_), .C(n951), .Y(n1172) );
  ao4f0 U1702 ( .A(n52), .B(n945), .C(n50), .D(n942), .Y(n1174) );
  ao4f0 U1703 ( .A(n53), .B(n934), .C(n54), .D(n933), .Y(n1176) );
  oa1d1 U1704 ( .A(n56), .B(n936), .C(n1176), .Y(n1177) );
  ao2i0 U1705 ( .A(n955), .B(alu_MuxB_11_), .C(n948), .D(n1178), .Y(n1179) );
  ao4f0 U1706 ( .A(n56), .B(n945), .C(n54), .D(n943), .Y(n1180) );
  ao4f0 U1707 ( .A(n57), .B(n934), .C(n58), .D(n932), .Y(n1182) );
  oa1d1 U1708 ( .A(n60), .B(n936), .C(n1182), .Y(n1183) );
  ao2i0 U1709 ( .A(n953), .B(alu_MuxB_12_), .C(n951), .D(n1184), .Y(n1185) );
  ao4f0 U1710 ( .A(n60), .B(n944), .C(n58), .D(n942), .Y(n1186) );
  ao4f0 U1711 ( .A(n61), .B(n934), .C(n62), .D(n1325), .Y(n1188) );
  oa1d1 U1712 ( .A(n64), .B(n936), .C(n1188), .Y(n1189) );
  ao2i0 U1713 ( .A(n954), .B(alu_MuxB_13_), .C(n950), .D(n1190), .Y(n1191) );
  ao4f0 U1714 ( .A(n64), .B(n945), .C(n62), .D(n942), .Y(n1192) );
  ao4f0 U1715 ( .A(n65), .B(n935), .C(n66), .D(n932), .Y(n1194) );
  oa1d1 U1716 ( .A(n68), .B(n936), .C(n1194), .Y(n1195) );
  ao2i0 U1717 ( .A(n952), .B(alu_MuxB_14_), .C(n950), .D(n1196), .Y(n1197) );
  ao4f0 U1718 ( .A(n68), .B(n944), .C(n66), .D(n943), .Y(n1198) );
  ao4f0 U1719 ( .A(n69), .B(n935), .C(n70), .D(n933), .Y(n1200) );
  oa1d1 U1720 ( .A(n72), .B(n1328), .C(n1200), .Y(n1201) );
  ao2i0 U1721 ( .A(n952), .B(alu_MuxB_15_), .C(n950), .D(n1202), .Y(n1203) );
  ao4f0 U1722 ( .A(n72), .B(n944), .C(n70), .D(n943), .Y(n1204) );
  ao4f0 U1723 ( .A(n73), .B(n934), .C(n74), .D(n933), .Y(n1206) );
  oa1d1 U1724 ( .A(n76), .B(n937), .C(n1206), .Y(n1207) );
  ao2i0 U1725 ( .A(n952), .B(alu_MuxB_16_), .C(n950), .D(n1208), .Y(n1209) );
  ao4f0 U1726 ( .A(n76), .B(n945), .C(n74), .D(n943), .Y(n1210) );
  ao4f0 U1727 ( .A(n77), .B(n935), .C(n78), .D(n1325), .Y(n1212) );
  oa1d1 U1728 ( .A(n80), .B(n936), .C(n1212), .Y(n1213) );
  ao2i0 U1729 ( .A(n952), .B(alu_MuxB_17_), .C(n950), .D(n1214), .Y(n1215) );
  ao4f0 U1730 ( .A(n80), .B(n944), .C(n78), .D(n943), .Y(n1216) );
  ao4f0 U1731 ( .A(n81), .B(n934), .C(n82), .D(n933), .Y(n1218) );
  oa1d1 U1732 ( .A(n84), .B(n1328), .C(n1218), .Y(n1219) );
  ao2i0 U1733 ( .A(n952), .B(alu_MuxB_18_), .C(n950), .D(n1220), .Y(n1221) );
  ao4f0 U1734 ( .A(n84), .B(n945), .C(n82), .D(n942), .Y(n1222) );
  ao4f0 U1735 ( .A(n85), .B(n935), .C(n86), .D(n933), .Y(n1224) );
  oa1d1 U1736 ( .A(n88), .B(n1328), .C(n1224), .Y(n1225) );
  ao2i0 U1737 ( .A(n952), .B(alu_MuxB_19_), .C(n950), .D(n1226), .Y(n1227) );
  ao4f0 U1738 ( .A(n12), .B(n944), .C(n10), .D(n942), .Y(n1228) );
  ao4f0 U1739 ( .A(n13), .B(n934), .C(n14), .D(n932), .Y(n1230) );
  oa1d1 U1740 ( .A(n16), .B(n1328), .C(n1230), .Y(n1231) );
  nand2a0 U1741 ( .A(n947), .B(alu_MuxB_1_), .Y(n1232) );
  ao2i0 U1742 ( .A(n952), .B(alu_MuxB_1_), .C(n950), .D(n1232), .Y(n1233) );
  ao4f0 U1743 ( .A(n88), .B(n945), .C(n86), .D(n942), .Y(n1234) );
  ao4f0 U1744 ( .A(n89), .B(n935), .C(n90), .D(n933), .Y(n1236) );
  oa1d1 U1745 ( .A(n92), .B(n1328), .C(n1236), .Y(n1237) );
  ao2i0 U1746 ( .A(n953), .B(alu_MuxB_20_), .C(n948), .D(n1238), .Y(n1239) );
  ao4f0 U1747 ( .A(n92), .B(n944), .C(n90), .D(n942), .Y(n1240) );
  ao4f0 U1748 ( .A(n93), .B(n934), .C(n94), .D(n932), .Y(n1242) );
  oa1d1 U1749 ( .A(n96), .B(n1328), .C(n1242), .Y(n1243) );
  ao2i0 U1750 ( .A(n953), .B(alu_MuxB_21_), .C(n950), .D(n1244), .Y(n1245) );
  ao4f0 U1751 ( .A(n96), .B(n944), .C(n94), .D(n942), .Y(n1246) );
  ao4f0 U1752 ( .A(n97), .B(n934), .C(n98), .D(n933), .Y(n1248) );
  oa1d1 U1753 ( .A(n100), .B(n1328), .C(n1248), .Y(n1249) );
  ao2i0 U1754 ( .A(n953), .B(alu_MuxB_22_), .C(n949), .D(n1250), .Y(n1251) );
  ao4f0 U1755 ( .A(n100), .B(n945), .C(n98), .D(n943), .Y(n1252) );
  ao4f0 U1756 ( .A(n101), .B(n935), .C(n102), .D(n932), .Y(n1254) );
  oa1d1 U1757 ( .A(n104), .B(n936), .C(n1254), .Y(n1255) );
  ao2i0 U1758 ( .A(n953), .B(alu_MuxB_23_), .C(n949), .D(n1256), .Y(n1257) );
  ao4f0 U1759 ( .A(n104), .B(n945), .C(n102), .D(n942), .Y(n1258) );
  ao4f0 U1760 ( .A(n105), .B(n1326), .C(n106), .D(n932), .Y(n1260) );
  oa1d1 U1761 ( .A(n108), .B(n937), .C(n1260), .Y(n1261) );
  ao2i0 U1762 ( .A(n953), .B(alu_MuxB_24_), .C(n1344), .D(n1262), .Y(n1263) );
  ao4f0 U1763 ( .A(n108), .B(n945), .C(n106), .D(n942), .Y(n1264) );
  ao4f0 U1764 ( .A(n109), .B(n935), .C(n110), .D(n933), .Y(n1266) );
  oa1d1 U1765 ( .A(n112), .B(n936), .C(n1266), .Y(n1267) );
  ao2i0 U1766 ( .A(n953), .B(alu_MuxB_25_), .C(n949), .D(n1268), .Y(n1269) );
  ao4f0 U1767 ( .A(n112), .B(n944), .C(n110), .D(n943), .Y(n1270) );
  ao2i0 U1768 ( .A(n954), .B(alu_MuxB_26_), .C(n949), .D(n1272), .Y(n1273) );
  ao4f0 U1769 ( .A(n124), .B(n945), .C(n122), .D(n942), .Y(n1274) );
  ao2i0 U1770 ( .A(n954), .B(alu_MuxB_27_), .C(n949), .D(n1276), .Y(n1277) );
  ao4f0 U1771 ( .A(n120), .B(n944), .C(n118), .D(n943), .Y(n1278) );
  ao2i0 U1772 ( .A(n954), .B(alu_MuxB_28_), .C(n949), .D(n1280), .Y(n1281) );
  ao4f0 U1773 ( .A(n116), .B(n944), .C(n114), .D(n1338), .Y(n1282) );
  ao2i0 U1774 ( .A(n954), .B(alu_MuxB_29_), .C(n949), .D(n1284), .Y(n1285) );
  ao4f0 U1775 ( .A(n16), .B(n944), .C(n14), .D(n942), .Y(n1286) );
  ao4f0 U1776 ( .A(n17), .B(n935), .C(n18), .D(n933), .Y(n1288) );
  oa1d1 U1777 ( .A(n20), .B(n937), .C(n1288), .Y(n1289) );
  nand2a0 U1778 ( .A(n946), .B(alu_MuxB_2_), .Y(n1290) );
  ao2i0 U1779 ( .A(n954), .B(alu_MuxB_2_), .C(n949), .D(n1290), .Y(n1291) );
  ao4f0 U1780 ( .A(n2), .B(n1338), .C(n4), .D(n945), .Y(n1292) );
  ao2i0 U1781 ( .A(n954), .B(alu_MuxB_30_), .C(n949), .D(n1294), .Y(n1295) );
  ao4f0 U1782 ( .A(n127), .B(n944), .C(n126), .D(n943), .Y(n1296) );
  mx2d0 U1783 ( .D0(n1298), .D1(n947), .S(alu_MuxB_31_), .Y(n1299) );
  ao4f0 U1784 ( .A(n20), .B(n944), .C(n18), .D(n1338), .Y(n1300) );
  ao4f0 U1785 ( .A(n21), .B(n1326), .C(n22), .D(n933), .Y(n1302) );
  oa1d1 U1786 ( .A(n24), .B(n936), .C(n1302), .Y(n1303) );
  ao2i0 U1787 ( .A(n954), .B(alu_MuxB_3_), .C(n949), .D(n1304), .Y(n1305) );
  ao4f0 U1788 ( .A(n24), .B(n944), .C(n22), .D(n943), .Y(n1306) );
  ao4f0 U1789 ( .A(n25), .B(n934), .C(n26), .D(n933), .Y(n1308) );
  oa1d1 U1790 ( .A(n28), .B(n936), .C(n1308), .Y(n1309) );
  ao2i0 U1791 ( .A(n955), .B(alu_MuxB_4_), .C(n949), .D(n1310), .Y(n1311) );
  ao4f0 U1792 ( .A(n28), .B(n945), .C(n26), .D(n943), .Y(n1312) );
  ao4f0 U1793 ( .A(n29), .B(n935), .C(n30), .D(n932), .Y(n1314) );
  oa1d1 U1794 ( .A(n32), .B(n937), .C(n1314), .Y(n1315) );
  ao4f0 U1795 ( .A(n32), .B(n945), .C(n30), .D(n943), .Y(n1316) );
  ao4f0 U1796 ( .A(n33), .B(n934), .C(n34), .D(n932), .Y(n1318) );
  oa1d1 U1797 ( .A(n36), .B(n1328), .C(n1318), .Y(n1319) );
  ao1f1 U1798 ( .A(n952), .B(alu_MuxA_6_), .C(n948), .Y(n1322) );
  ao2i0 U1799 ( .A(n955), .B(alu_MuxB_6_), .C(n949), .D(n1320), .Y(n1321) );
  ao4f0 U1800 ( .A(n36), .B(n944), .C(n34), .D(n943), .Y(n1323) );
  ao4f0 U1801 ( .A(n37), .B(n935), .C(n38), .D(n933), .Y(n1327) );
  oa1d1 U1802 ( .A(n40), .B(n1328), .C(n1327), .Y(n1329) );
  ao2i0 U1803 ( .A(n955), .B(alu_MuxB_7_), .C(n951), .D(n1331), .Y(n1332) );
  ao4f0 U1804 ( .A(n40), .B(n1339), .C(n38), .D(n942), .Y(n1333) );
  ao2i0 U1805 ( .A(n955), .B(alu_MuxB_8_), .C(n1344), .D(n1335), .Y(n1336) );
  ao4f0 U1806 ( .A(n44), .B(n945), .C(n42), .D(n943), .Y(n1340) );
  ao2i0 U1807 ( .A(n952), .B(alu_MuxB_9_), .C(n949), .D(n1343), .Y(n1346) );
  oa2i0 U1808 ( .A(cntrl_state_2_), .B(n419), .C(cntrl_state_7_), .D(n426), 
        .Y(n1348) );
  oa1d1 U1809 ( .A(cntrl_state_9_), .B(cntrl_state_8_), .C(Reset), .Y(
        cntrl_N111) );
  mx2d0 U1810 ( .D0(n1481), .D1(n128), .S(n963), .Y(n895) );
  and3d1 U1811 ( .A(n1437), .B(PCSource[0]), .C(PCSource[1]), .Y(n1439) );
  oa4f0 U1812 ( .A(PC[1]), .B(n958), .C(n959), .D(TargetReg[1]), .Y(n1379) );
  ao2i0 U1813 ( .A(n957), .B(n1148), .C(n1379), .D(n1378), .Y(n893) );
  oa4f0 U1814 ( .A(PC[2]), .B(n1437), .C(n1438), .D(TargetReg[2]), .Y(n1381)
         );
  nand2a0 U1815 ( .A(n960), .B(WriteAdd[2]), .Y(n1380) );
  ao2i0 U1816 ( .A(n957), .B(n1149), .C(n1381), .D(n1380), .Y(n892) );
  oa4f0 U1817 ( .A(Instruction[3]), .B(n956), .C(PC[3]), .D(n958), .Y(n1383)
         );
  oa4f0 U1818 ( .A(TargetReg[3]), .B(n1438), .C(n960), .D(WriteAdd[3]), .Y(
        n1382) );
  oa4f0 U1819 ( .A(Instruction[4]), .B(n956), .C(PC[4]), .D(n958), .Y(n1385)
         );
  oa4f0 U1820 ( .A(TargetReg[4]), .B(n959), .C(n960), .D(WriteAdd[4]), .Y(
        n1384) );
  oa4f0 U1821 ( .A(Instruction[5]), .B(n1434), .C(PC[5]), .D(n958), .Y(n1387)
         );
  oa4f0 U1822 ( .A(TargetReg[5]), .B(n1438), .C(n960), .D(WriteAdd[5]), .Y(
        n1386) );
  oa4f0 U1823 ( .A(Instruction[6]), .B(n1434), .C(PC[6]), .D(n958), .Y(n1389)
         );
  oa4f0 U1824 ( .A(TargetReg[6]), .B(n959), .C(n960), .D(WriteAdd[6]), .Y(
        n1388) );
  oa4f0 U1825 ( .A(Instruction[7]), .B(n1434), .C(PC[7]), .D(n958), .Y(n1391)
         );
  oa4f0 U1826 ( .A(TargetReg[7]), .B(n959), .C(n960), .D(WriteAdd[7]), .Y(
        n1390) );
  oa4f0 U1827 ( .A(Instruction[8]), .B(n1434), .C(PC[8]), .D(n958), .Y(n1393)
         );
  oa4f0 U1828 ( .A(TargetReg[8]), .B(n959), .C(n960), .D(WriteAdd[8]), .Y(
        n1392) );
  oa4f0 U1829 ( .A(Instruction[9]), .B(n1434), .C(PC[9]), .D(n1437), .Y(n1395)
         );
  oa4f0 U1830 ( .A(TargetReg[9]), .B(n959), .C(n1439), .D(WriteAdd[9]), .Y(
        n1394) );
  oa4f0 U1831 ( .A(Instruction[10]), .B(n1434), .C(PC[10]), .D(n958), .Y(n1397) );
  oa4f0 U1832 ( .A(TargetReg[10]), .B(n1438), .C(n960), .D(WriteAdd[10]), .Y(
        n1396) );
  oa4f0 U1833 ( .A(Instruction[11]), .B(n1434), .C(PC[11]), .D(n958), .Y(n1399) );
  oa4f0 U1834 ( .A(TargetReg[11]), .B(n959), .C(n960), .D(WriteAdd[11]), .Y(
        n1398) );
  oa4f0 U1835 ( .A(Instruction[12]), .B(n1434), .C(PC[12]), .D(n958), .Y(n1401) );
  oa4f0 U1836 ( .A(TargetReg[12]), .B(n1438), .C(n1439), .D(WriteAdd[12]), .Y(
        n1400) );
  oa4f0 U1837 ( .A(Instruction[13]), .B(n1434), .C(PC[13]), .D(n1437), .Y(
        n1403) );
  oa4f0 U1838 ( .A(TargetReg[13]), .B(n959), .C(n960), .D(WriteAdd[13]), .Y(
        n1402) );
  oa4f0 U1839 ( .A(Instruction[14]), .B(n1434), .C(PC[14]), .D(n958), .Y(n1405) );
  oa4f0 U1840 ( .A(TargetReg[14]), .B(n1438), .C(n1439), .D(WriteAdd[14]), .Y(
        n1404) );
  oa4f0 U1841 ( .A(Instruction[15]), .B(n956), .C(PC[15]), .D(n958), .Y(n1407)
         );
  oa4f0 U1842 ( .A(TargetReg[15]), .B(n1438), .C(n1439), .D(WriteAdd[15]), .Y(
        n1406) );
  oa4f0 U1843 ( .A(Read2RegSel[0]), .B(n956), .C(PC[16]), .D(n1437), .Y(n1409)
         );
  oa4f0 U1844 ( .A(TargetReg[16]), .B(n959), .C(n960), .D(WriteAdd[16]), .Y(
        n1408) );
  oa4f0 U1845 ( .A(Read2RegSel[1]), .B(n956), .C(PC[17]), .D(n958), .Y(n1411)
         );
  oa4f0 U1846 ( .A(TargetReg[17]), .B(n959), .C(n960), .D(WriteAdd[17]), .Y(
        n1410) );
  oa4f0 U1847 ( .A(PC[18]), .B(n1437), .C(n1434), .D(Instruction_18), .Y(n1413) );
  oa4f0 U1848 ( .A(TargetReg[18]), .B(n1438), .C(n960), .D(WriteAdd[18]), .Y(
        n1412) );
  oa4f0 U1849 ( .A(PC[19]), .B(n958), .C(n956), .D(Instruction_19), .Y(n1415)
         );
  oa4f0 U1850 ( .A(TargetReg[19]), .B(n1438), .C(n960), .D(WriteAdd[19]), .Y(
        n1414) );
  oa4f0 U1851 ( .A(PC[20]), .B(n958), .C(n1434), .D(Instruction_20), .Y(n1417)
         );
  oa4f0 U1852 ( .A(TargetReg[20]), .B(n959), .C(n1439), .D(WriteAdd[20]), .Y(
        n1416) );
  oa4f0 U1853 ( .A(Read1RegSel[0]), .B(n1434), .C(PC[21]), .D(n958), .Y(n1419)
         );
  oa4f0 U1854 ( .A(TargetReg[21]), .B(n959), .C(n1439), .D(WriteAdd[21]), .Y(
        n1418) );
  oa4f0 U1855 ( .A(Read1RegSel[1]), .B(n1434), .C(PC[22]), .D(n958), .Y(n1421)
         );
  oa4f0 U1856 ( .A(TargetReg[22]), .B(n959), .C(n960), .D(WriteAdd[22]), .Y(
        n1420) );
  oa4f0 U1857 ( .A(PC[23]), .B(n1437), .C(n956), .D(Instruction_23), .Y(n1423)
         );
  oa4f0 U1858 ( .A(TargetReg[23]), .B(n959), .C(n1439), .D(WriteAdd[23]), .Y(
        n1422) );
  oa4f0 U1859 ( .A(PC[24]), .B(n1437), .C(n956), .D(Instruction_24), .Y(n1425)
         );
  oa4f0 U1860 ( .A(TargetReg[24]), .B(n1438), .C(n960), .D(WriteAdd[24]), .Y(
        n1424) );
  oa4f0 U1861 ( .A(PC[25]), .B(n1437), .C(n956), .D(Instruction_25), .Y(n1427)
         );
  oa4f0 U1862 ( .A(TargetReg[25]), .B(n1438), .C(n960), .D(WriteAdd[25]), .Y(
        n1426) );
  oa4f0 U1863 ( .A(PC[28]), .B(n1434), .C(PC[26]), .D(n958), .Y(n1429) );
  oa4f0 U1864 ( .A(TargetReg[26]), .B(n1438), .C(n960), .D(WriteAdd[26]), .Y(
        n1428) );
  oa4f0 U1865 ( .A(PC[29]), .B(n956), .C(PC[27]), .D(n958), .Y(n1431) );
  oa4f0 U1866 ( .A(TargetReg[27]), .B(n1438), .C(n960), .D(WriteAdd[27]), .Y(
        n1430) );
  oa4f0 U1867 ( .A(PC[30]), .B(n956), .C(PC[28]), .D(n958), .Y(n1433) );
  oa4f0 U1868 ( .A(TargetReg[28]), .B(n959), .C(n960), .D(WriteAdd[28]), .Y(
        n1432) );
  oa4f0 U1869 ( .A(PC[29]), .B(n1437), .C(PC[31]), .D(n1434), .Y(n1436) );
  oa4f0 U1870 ( .A(TargetReg[29]), .B(n1438), .C(n1439), .D(WriteAdd[29]), .Y(
        n1435) );
  mx2d0 U1871 ( .D0(n1445), .D1(n5), .S(n965), .Y(n862) );
  mx2d0 U1872 ( .D0(n1445), .D1(n6), .S(n968), .Y(n861) );
  mx2d0 U1873 ( .D0(n1445), .D1(n7), .S(n964), .Y(n860) );
  mx2d0 U1874 ( .D0(n1445), .D1(n8), .S(n970), .Y(n859) );
  mx2d0 U1875 ( .D0(n1446), .D1(n9), .S(n966), .Y(n858) );
  mx2d0 U1876 ( .D0(n1446), .D1(n10), .S(n967), .Y(n857) );
  mx2d0 U1877 ( .D0(n1446), .D1(n11), .S(n963), .Y(n856) );
  mx2d0 U1878 ( .D0(n1446), .D1(n12), .S(n969), .Y(n855) );
  mx2d0 U1879 ( .D0(n1447), .D1(n13), .S(n965), .Y(n854) );
  mx2d0 U1880 ( .D0(n1447), .D1(n14), .S(n968), .Y(n853) );
  mx2d0 U1881 ( .D0(n1447), .D1(n15), .S(n963), .Y(n852) );
  mx2d0 U1882 ( .D0(n1447), .D1(n16), .S(n970), .Y(n851) );
  mx2d0 U1883 ( .D0(n1448), .D1(n17), .S(n965), .Y(n850) );
  mx2d0 U1884 ( .D0(n1448), .D1(n18), .S(n968), .Y(n849) );
  mx2d0 U1885 ( .D0(n1448), .D1(n19), .S(n963), .Y(n848) );
  mx2d0 U1886 ( .D0(n1448), .D1(n20), .S(n970), .Y(n847) );
  mx2d0 U1887 ( .D0(n1449), .D1(n21), .S(n965), .Y(n846) );
  mx2d0 U1888 ( .D0(n1449), .D1(n22), .S(n968), .Y(n845) );
  mx2d0 U1889 ( .D0(n1449), .D1(n23), .S(n963), .Y(n844) );
  mx2d0 U1890 ( .D0(n1449), .D1(n24), .S(n970), .Y(n843) );
  mx2d0 U1891 ( .D0(n1450), .D1(n25), .S(n965), .Y(n842) );
  mx2d0 U1892 ( .D0(n1450), .D1(n26), .S(n1479), .Y(n841) );
  mx2d0 U1893 ( .D0(n1450), .D1(n27), .S(n964), .Y(n840) );
  mx2d0 U1894 ( .D0(n1450), .D1(n28), .S(n1480), .Y(n839) );
  mx2d0 U1895 ( .D0(n1451), .D1(n29), .S(n966), .Y(n838) );
  mx2d0 U1896 ( .D0(n1451), .D1(n30), .S(n967), .Y(n837) );
  mx2d0 U1897 ( .D0(n1451), .D1(n31), .S(n963), .Y(n836) );
  mx2d0 U1898 ( .D0(n1451), .D1(n32), .S(n969), .Y(n835) );
  mx2d0 U1899 ( .D0(n1452), .D1(n33), .S(n965), .Y(n834) );
  mx2d0 U1900 ( .D0(n1452), .D1(n34), .S(n967), .Y(n833) );
  mx2d0 U1901 ( .D0(n1452), .D1(n35), .S(n1476), .Y(n832) );
  mx2d0 U1902 ( .D0(n1452), .D1(n36), .S(n969), .Y(n831) );
  mx2d0 U1903 ( .D0(n1453), .D1(n37), .S(n1478), .Y(n830) );
  mx2d0 U1904 ( .D0(n1453), .D1(n38), .S(n968), .Y(n829) );
  mx2d0 U1905 ( .D0(n1453), .D1(n39), .S(n964), .Y(n828) );
  mx2d0 U1906 ( .D0(n1453), .D1(n40), .S(n970), .Y(n827) );
  mx2d0 U1907 ( .D0(n1454), .D1(n41), .S(n966), .Y(n826) );
  mx2d0 U1908 ( .D0(n1454), .D1(n42), .S(n968), .Y(n825) );
  mx2d0 U1909 ( .D0(n1454), .D1(n43), .S(n963), .Y(n824) );
  mx2d0 U1910 ( .D0(n1454), .D1(n44), .S(n970), .Y(n823) );
  mx2d0 U1911 ( .D0(n1455), .D1(n45), .S(n965), .Y(n822) );
  mx2d0 U1912 ( .D0(n1455), .D1(n47), .S(n963), .Y(n820) );
  mx2d0 U1913 ( .D0(n1456), .D1(n49), .S(n965), .Y(n818) );
  mx2d0 U1914 ( .D0(n1456), .D1(n50), .S(n968), .Y(n817) );
  mx2d0 U1915 ( .D0(n1456), .D1(n51), .S(n964), .Y(n816) );
  mx2d0 U1916 ( .D0(n1456), .D1(n52), .S(n970), .Y(n815) );
  mx2d0 U1917 ( .D0(n1457), .D1(n53), .S(n966), .Y(n814) );
  mx2d0 U1918 ( .D0(n1457), .D1(n54), .S(n967), .Y(n813) );
  mx2d0 U1919 ( .D0(n1457), .D1(n55), .S(n964), .Y(n812) );
  mx2d0 U1920 ( .D0(n1457), .D1(n56), .S(n969), .Y(n811) );
  mx2d0 U1921 ( .D0(n1458), .D1(n57), .S(n966), .Y(n810) );
  mx2d0 U1922 ( .D0(n1458), .D1(n58), .S(n967), .Y(n809) );
  mx2d0 U1923 ( .D0(n1458), .D1(n59), .S(n964), .Y(n808) );
  mx2d0 U1924 ( .D0(n1458), .D1(n60), .S(n969), .Y(n807) );
  mx2d0 U1925 ( .D0(n1459), .D1(n61), .S(n966), .Y(n806) );
  mx2d0 U1926 ( .D0(n1459), .D1(n62), .S(n967), .Y(n805) );
  mx2d0 U1927 ( .D0(n1459), .D1(n63), .S(n964), .Y(n804) );
  mx2d0 U1928 ( .D0(n1459), .D1(n64), .S(n969), .Y(n803) );
  mx2d0 U1929 ( .D0(n1460), .D1(n65), .S(n966), .Y(n802) );
  mx2d0 U1930 ( .D0(n1460), .D1(n66), .S(n967), .Y(n801) );
  mx2d0 U1931 ( .D0(n1460), .D1(n67), .S(n964), .Y(n800) );
  mx2d0 U1932 ( .D0(n1460), .D1(n68), .S(n969), .Y(n799) );
  mx2d0 U1933 ( .D0(n1461), .D1(n69), .S(n966), .Y(n798) );
  mx2d0 U1934 ( .D0(n1461), .D1(n70), .S(n967), .Y(n797) );
  mx2d0 U1935 ( .D0(n1461), .D1(n71), .S(n964), .Y(n796) );
  mx2d0 U1936 ( .D0(n1461), .D1(n72), .S(n969), .Y(n795) );
  mx2d0 U1937 ( .D0(n1462), .D1(n73), .S(n966), .Y(n794) );
  mx2d0 U1938 ( .D0(n1462), .D1(n74), .S(n967), .Y(n793) );
  mx2d0 U1939 ( .D0(n1462), .D1(n75), .S(n1476), .Y(n792) );
  mx2d0 U1940 ( .D0(n1462), .D1(n76), .S(n969), .Y(n791) );
  mx2d0 U1941 ( .D0(n1463), .D1(n77), .S(n1478), .Y(n790) );
  mx2d0 U1942 ( .D0(n1463), .D1(n78), .S(n967), .Y(n789) );
  mx2d0 U1943 ( .D0(n1463), .D1(n79), .S(n963), .Y(n788) );
  mx2d0 U1944 ( .D0(n1463), .D1(n80), .S(n969), .Y(n787) );
  mx2d0 U1945 ( .D0(n1464), .D1(n81), .S(n965), .Y(n786) );
  mx2d0 U1946 ( .D0(n1464), .D1(n82), .S(n968), .Y(n785) );
  mx2d0 U1947 ( .D0(n1464), .D1(n83), .S(n1476), .Y(n784) );
  mx2d0 U1948 ( .D0(n1464), .D1(n84), .S(n970), .Y(n783) );
  mx2d0 U1949 ( .D0(n1465), .D1(n85), .S(n1478), .Y(n782) );
  mx2d0 U1950 ( .D0(n1465), .D1(n86), .S(n1479), .Y(n781) );
  mx2d0 U1951 ( .D0(n1465), .D1(n87), .S(n1476), .Y(n780) );
  mx2d0 U1952 ( .D0(n1465), .D1(n88), .S(n1480), .Y(n779) );
  mx2d0 U1953 ( .D0(n1466), .D1(n89), .S(n1478), .Y(n778) );
  mx2d0 U1954 ( .D0(n1466), .D1(n90), .S(n1479), .Y(n777) );
  mx2d0 U1955 ( .D0(n1466), .D1(n91), .S(n964), .Y(n776) );
  mx2d0 U1956 ( .D0(n1466), .D1(n92), .S(n1480), .Y(n775) );
  mx2d0 U1957 ( .D0(n1467), .D1(n93), .S(n966), .Y(n774) );
  mx2d0 U1958 ( .D0(n1467), .D1(n94), .S(n1479), .Y(n773) );
  mx2d0 U1959 ( .D0(n1467), .D1(n95), .S(n963), .Y(n772) );
  mx2d0 U1960 ( .D0(n1467), .D1(n96), .S(n1480), .Y(n771) );
  mx2d0 U1961 ( .D0(n1468), .D1(n97), .S(n965), .Y(n770) );
  mx2d0 U1962 ( .D0(n1468), .D1(n98), .S(n1479), .Y(n769) );
  mx2d0 U1963 ( .D0(n1468), .D1(n99), .S(n1476), .Y(n768) );
  mx2d0 U1964 ( .D0(n1468), .D1(n100), .S(n1480), .Y(n767) );
  mx2d0 U1965 ( .D0(n1469), .D1(n101), .S(n1478), .Y(n766) );
  mx2d0 U1966 ( .D0(n1469), .D1(n102), .S(n968), .Y(n765) );
  mx2d0 U1967 ( .D0(n1469), .D1(n103), .S(n964), .Y(n764) );
  mx2d0 U1968 ( .D0(n1469), .D1(n104), .S(n970), .Y(n763) );
  mx2d0 U1969 ( .D0(n1470), .D1(n105), .S(n966), .Y(n762) );
  mx2d0 U1970 ( .D0(n1470), .D1(n106), .S(n967), .Y(n761) );
  mx2d0 U1971 ( .D0(n1470), .D1(n107), .S(n963), .Y(n760) );
  mx2d0 U1972 ( .D0(n1470), .D1(n108), .S(n969), .Y(n759) );
  mx2d0 U1973 ( .D0(n1471), .D1(n109), .S(n965), .Y(n758) );
  mx2d0 U1974 ( .D0(n1471), .D1(n110), .S(n968), .Y(n757) );
  mx2d0 U1975 ( .D0(n1471), .D1(n111), .S(n1476), .Y(n756) );
  mx2d0 U1976 ( .D0(n1471), .D1(n112), .S(n970), .Y(n755) );
  mx2d0 U1977 ( .D0(n1472), .D1(n121), .S(n1478), .Y(n754) );
  mx2d0 U1978 ( .D0(n1472), .D1(n122), .S(n1479), .Y(n753) );
  mx2d0 U1979 ( .D0(n1472), .D1(n123), .S(n964), .Y(n752) );
  mx2d0 U1980 ( .D0(n1472), .D1(n124), .S(n1480), .Y(n751) );
  mx2d0 U1981 ( .D0(n1473), .D1(n117), .S(n966), .Y(n750) );
  mx2d0 U1982 ( .D0(n1473), .D1(n118), .S(n967), .Y(n749) );
  mx2d0 U1983 ( .D0(n1473), .D1(n119), .S(n963), .Y(n748) );
  mx2d0 U1984 ( .D0(n1473), .D1(n120), .S(n969), .Y(n747) );
  mx2d0 U1985 ( .D0(n1474), .D1(n113), .S(n965), .Y(n746) );
  mx2d0 U1986 ( .D0(n1474), .D1(n114), .S(n968), .Y(n745) );
  mx2d0 U1987 ( .D0(n1474), .D1(n115), .S(n1476), .Y(n744) );
  mx2d0 U1988 ( .D0(n1474), .D1(n116), .S(n970), .Y(n743) );
  mx2d0 U1989 ( .D0(n1477), .D1(n1), .S(n1478), .Y(n742) );
  mx2d0 U1990 ( .D0(n1477), .D1(n2), .S(n1479), .Y(n741) );
  mx2d0 U1991 ( .D0(n1477), .D1(n3), .S(n1476), .Y(n740) );
  mx2d0 U1992 ( .D0(n1477), .D1(n4), .S(n1480), .Y(n739) );
  mx2d0 U1993 ( .D0(n1481), .D1(n125), .S(n1478), .Y(n738) );
  mx2d0 U1994 ( .D0(n1481), .D1(n126), .S(n1479), .Y(n737) );
  mx2d0 U1995 ( .D0(n1481), .D1(n127), .S(n1480), .Y(n736) );
endmodule

